
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c4",x"f2",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c4",x"f2",x"c2"),
    14 => (x"48",x"cc",x"df",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"d9",x"e2"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"c4",x"4a",x"71",x"1e"),
    47 => (x"c1",x"48",x"49",x"66"),
    48 => (x"58",x"a6",x"c8",x"88"),
    49 => (x"d4",x"02",x"99",x"71"),
    50 => (x"ff",x"48",x"12",x"87"),
    51 => (x"c4",x"78",x"08",x"d4"),
    52 => (x"c1",x"48",x"49",x"66"),
    53 => (x"58",x"a6",x"c8",x"88"),
    54 => (x"ec",x"05",x"99",x"71"),
    55 => (x"1e",x"4f",x"26",x"87"),
    56 => (x"66",x"c4",x"4a",x"71"),
    57 => (x"88",x"c1",x"48",x"49"),
    58 => (x"71",x"58",x"a6",x"c8"),
    59 => (x"87",x"d6",x"02",x"99"),
    60 => (x"c3",x"48",x"d4",x"ff"),
    61 => (x"52",x"68",x"78",x"ff"),
    62 => (x"48",x"49",x"66",x"c4"),
    63 => (x"a6",x"c8",x"88",x"c1"),
    64 => (x"05",x"99",x"71",x"58"),
    65 => (x"4f",x"26",x"87",x"ea"),
    66 => (x"ff",x"1e",x"73",x"1e"),
    67 => (x"ff",x"c3",x"4b",x"d4"),
    68 => (x"c3",x"4a",x"6b",x"7b"),
    69 => (x"49",x"6b",x"7b",x"ff"),
    70 => (x"b1",x"72",x"32",x"c8"),
    71 => (x"6b",x"7b",x"ff",x"c3"),
    72 => (x"71",x"31",x"c8",x"4a"),
    73 => (x"7b",x"ff",x"c3",x"b2"),
    74 => (x"32",x"c8",x"49",x"6b"),
    75 => (x"48",x"71",x"b1",x"72"),
    76 => (x"4d",x"26",x"87",x"c4"),
    77 => (x"4b",x"26",x"4c",x"26"),
    78 => (x"5e",x"0e",x"4f",x"26"),
    79 => (x"0e",x"5d",x"5c",x"5b"),
    80 => (x"d4",x"ff",x"4a",x"71"),
    81 => (x"c3",x"49",x"72",x"4c"),
    82 => (x"7c",x"71",x"99",x"ff"),
    83 => (x"bf",x"cc",x"df",x"c2"),
    84 => (x"d0",x"87",x"c8",x"05"),
    85 => (x"30",x"c9",x"48",x"66"),
    86 => (x"d0",x"58",x"a6",x"d4"),
    87 => (x"29",x"d8",x"49",x"66"),
    88 => (x"71",x"99",x"ff",x"c3"),
    89 => (x"49",x"66",x"d0",x"7c"),
    90 => (x"ff",x"c3",x"29",x"d0"),
    91 => (x"d0",x"7c",x"71",x"99"),
    92 => (x"29",x"c8",x"49",x"66"),
    93 => (x"71",x"99",x"ff",x"c3"),
    94 => (x"49",x"66",x"d0",x"7c"),
    95 => (x"71",x"99",x"ff",x"c3"),
    96 => (x"d0",x"49",x"72",x"7c"),
    97 => (x"99",x"ff",x"c3",x"29"),
    98 => (x"4b",x"6c",x"7c",x"71"),
    99 => (x"4d",x"ff",x"f0",x"c9"),
   100 => (x"05",x"ab",x"ff",x"c3"),
   101 => (x"ff",x"c3",x"87",x"d0"),
   102 => (x"c1",x"4b",x"6c",x"7c"),
   103 => (x"87",x"c6",x"02",x"8d"),
   104 => (x"02",x"ab",x"ff",x"c3"),
   105 => (x"48",x"73",x"87",x"f0"),
   106 => (x"1e",x"87",x"c7",x"fe"),
   107 => (x"d4",x"ff",x"49",x"c0"),
   108 => (x"78",x"ff",x"c3",x"48"),
   109 => (x"c8",x"c3",x"81",x"c1"),
   110 => (x"f1",x"04",x"a9",x"b7"),
   111 => (x"1e",x"4f",x"26",x"87"),
   112 => (x"87",x"e7",x"1e",x"73"),
   113 => (x"4b",x"df",x"f8",x"c4"),
   114 => (x"ff",x"c0",x"1e",x"c0"),
   115 => (x"49",x"f7",x"c1",x"f0"),
   116 => (x"c4",x"87",x"e7",x"fd"),
   117 => (x"05",x"a8",x"c1",x"86"),
   118 => (x"ff",x"87",x"ea",x"c0"),
   119 => (x"ff",x"c3",x"48",x"d4"),
   120 => (x"c0",x"c0",x"c1",x"78"),
   121 => (x"1e",x"c0",x"c0",x"c0"),
   122 => (x"c1",x"f0",x"e1",x"c0"),
   123 => (x"c9",x"fd",x"49",x"e9"),
   124 => (x"70",x"86",x"c4",x"87"),
   125 => (x"87",x"ca",x"05",x"98"),
   126 => (x"c3",x"48",x"d4",x"ff"),
   127 => (x"48",x"c1",x"78",x"ff"),
   128 => (x"e6",x"fe",x"87",x"cb"),
   129 => (x"05",x"8b",x"c1",x"87"),
   130 => (x"c0",x"87",x"fd",x"fe"),
   131 => (x"87",x"e6",x"fc",x"48"),
   132 => (x"ff",x"1e",x"73",x"1e"),
   133 => (x"ff",x"c3",x"48",x"d4"),
   134 => (x"c0",x"4b",x"d3",x"78"),
   135 => (x"f0",x"ff",x"c0",x"1e"),
   136 => (x"fc",x"49",x"c1",x"c1"),
   137 => (x"86",x"c4",x"87",x"d4"),
   138 => (x"ca",x"05",x"98",x"70"),
   139 => (x"48",x"d4",x"ff",x"87"),
   140 => (x"c1",x"78",x"ff",x"c3"),
   141 => (x"fd",x"87",x"cb",x"48"),
   142 => (x"8b",x"c1",x"87",x"f1"),
   143 => (x"87",x"db",x"ff",x"05"),
   144 => (x"f1",x"fb",x"48",x"c0"),
   145 => (x"5b",x"5e",x"0e",x"87"),
   146 => (x"d4",x"ff",x"0e",x"5c"),
   147 => (x"87",x"db",x"fd",x"4c"),
   148 => (x"c0",x"1e",x"ea",x"c6"),
   149 => (x"c8",x"c1",x"f0",x"e1"),
   150 => (x"87",x"de",x"fb",x"49"),
   151 => (x"a8",x"c1",x"86",x"c4"),
   152 => (x"fe",x"87",x"c8",x"02"),
   153 => (x"48",x"c0",x"87",x"ea"),
   154 => (x"fa",x"87",x"e2",x"c1"),
   155 => (x"49",x"70",x"87",x"da"),
   156 => (x"99",x"ff",x"ff",x"cf"),
   157 => (x"02",x"a9",x"ea",x"c6"),
   158 => (x"d3",x"fe",x"87",x"c8"),
   159 => (x"c1",x"48",x"c0",x"87"),
   160 => (x"ff",x"c3",x"87",x"cb"),
   161 => (x"4b",x"f1",x"c0",x"7c"),
   162 => (x"70",x"87",x"f4",x"fc"),
   163 => (x"eb",x"c0",x"02",x"98"),
   164 => (x"c0",x"1e",x"c0",x"87"),
   165 => (x"fa",x"c1",x"f0",x"ff"),
   166 => (x"87",x"de",x"fa",x"49"),
   167 => (x"98",x"70",x"86",x"c4"),
   168 => (x"c3",x"87",x"d9",x"05"),
   169 => (x"49",x"6c",x"7c",x"ff"),
   170 => (x"7c",x"7c",x"ff",x"c3"),
   171 => (x"c0",x"c1",x"7c",x"7c"),
   172 => (x"87",x"c4",x"02",x"99"),
   173 => (x"87",x"d5",x"48",x"c1"),
   174 => (x"87",x"d1",x"48",x"c0"),
   175 => (x"c4",x"05",x"ab",x"c2"),
   176 => (x"c8",x"48",x"c0",x"87"),
   177 => (x"05",x"8b",x"c1",x"87"),
   178 => (x"c0",x"87",x"fd",x"fe"),
   179 => (x"87",x"e4",x"f9",x"48"),
   180 => (x"c2",x"1e",x"73",x"1e"),
   181 => (x"c1",x"48",x"cc",x"df"),
   182 => (x"ff",x"4b",x"c7",x"78"),
   183 => (x"78",x"c2",x"48",x"d0"),
   184 => (x"ff",x"87",x"c8",x"fb"),
   185 => (x"78",x"c3",x"48",x"d0"),
   186 => (x"e5",x"c0",x"1e",x"c0"),
   187 => (x"49",x"c0",x"c1",x"d0"),
   188 => (x"c4",x"87",x"c7",x"f9"),
   189 => (x"05",x"a8",x"c1",x"86"),
   190 => (x"c2",x"4b",x"87",x"c1"),
   191 => (x"87",x"c5",x"05",x"ab"),
   192 => (x"f9",x"c0",x"48",x"c0"),
   193 => (x"05",x"8b",x"c1",x"87"),
   194 => (x"fc",x"87",x"d0",x"ff"),
   195 => (x"df",x"c2",x"87",x"f7"),
   196 => (x"98",x"70",x"58",x"d0"),
   197 => (x"c1",x"87",x"cd",x"05"),
   198 => (x"f0",x"ff",x"c0",x"1e"),
   199 => (x"f8",x"49",x"d0",x"c1"),
   200 => (x"86",x"c4",x"87",x"d8"),
   201 => (x"c3",x"48",x"d4",x"ff"),
   202 => (x"de",x"c4",x"78",x"ff"),
   203 => (x"d4",x"df",x"c2",x"87"),
   204 => (x"48",x"d0",x"ff",x"58"),
   205 => (x"d4",x"ff",x"78",x"c2"),
   206 => (x"78",x"ff",x"c3",x"48"),
   207 => (x"f5",x"f7",x"48",x"c1"),
   208 => (x"5b",x"5e",x"0e",x"87"),
   209 => (x"71",x"0e",x"5d",x"5c"),
   210 => (x"4d",x"ff",x"c3",x"4a"),
   211 => (x"75",x"4c",x"d4",x"ff"),
   212 => (x"48",x"d0",x"ff",x"7c"),
   213 => (x"75",x"78",x"c3",x"c4"),
   214 => (x"c0",x"1e",x"72",x"7c"),
   215 => (x"d8",x"c1",x"f0",x"ff"),
   216 => (x"87",x"d6",x"f7",x"49"),
   217 => (x"98",x"70",x"86",x"c4"),
   218 => (x"c1",x"87",x"c5",x"02"),
   219 => (x"87",x"f0",x"c0",x"48"),
   220 => (x"fe",x"c3",x"7c",x"75"),
   221 => (x"1e",x"c0",x"c8",x"7c"),
   222 => (x"f4",x"49",x"66",x"d4"),
   223 => (x"86",x"c4",x"87",x"fa"),
   224 => (x"7c",x"75",x"7c",x"75"),
   225 => (x"da",x"d8",x"7c",x"75"),
   226 => (x"7c",x"75",x"4b",x"e0"),
   227 => (x"05",x"99",x"49",x"6c"),
   228 => (x"8b",x"c1",x"87",x"c5"),
   229 => (x"75",x"87",x"f3",x"05"),
   230 => (x"48",x"d0",x"ff",x"7c"),
   231 => (x"48",x"c0",x"78",x"c2"),
   232 => (x"0e",x"87",x"cf",x"f6"),
   233 => (x"5d",x"5c",x"5b",x"5e"),
   234 => (x"c0",x"4b",x"71",x"0e"),
   235 => (x"cd",x"ee",x"c5",x"4c"),
   236 => (x"d4",x"ff",x"4a",x"df"),
   237 => (x"78",x"ff",x"c3",x"48"),
   238 => (x"fe",x"c3",x"49",x"68"),
   239 => (x"fd",x"c0",x"05",x"a9"),
   240 => (x"73",x"4d",x"70",x"87"),
   241 => (x"87",x"cc",x"02",x"9b"),
   242 => (x"73",x"1e",x"66",x"d0"),
   243 => (x"87",x"cf",x"f4",x"49"),
   244 => (x"87",x"d6",x"86",x"c4"),
   245 => (x"c4",x"48",x"d0",x"ff"),
   246 => (x"ff",x"c3",x"78",x"d1"),
   247 => (x"48",x"66",x"d0",x"7d"),
   248 => (x"a6",x"d4",x"88",x"c1"),
   249 => (x"05",x"98",x"70",x"58"),
   250 => (x"d4",x"ff",x"87",x"f0"),
   251 => (x"78",x"ff",x"c3",x"48"),
   252 => (x"05",x"9b",x"73",x"78"),
   253 => (x"d0",x"ff",x"87",x"c5"),
   254 => (x"c1",x"78",x"d0",x"48"),
   255 => (x"8a",x"c1",x"4c",x"4a"),
   256 => (x"87",x"ee",x"fe",x"05"),
   257 => (x"e9",x"f4",x"48",x"74"),
   258 => (x"1e",x"73",x"1e",x"87"),
   259 => (x"4b",x"c0",x"4a",x"71"),
   260 => (x"c3",x"48",x"d4",x"ff"),
   261 => (x"d0",x"ff",x"78",x"ff"),
   262 => (x"78",x"c3",x"c4",x"48"),
   263 => (x"c3",x"48",x"d4",x"ff"),
   264 => (x"1e",x"72",x"78",x"ff"),
   265 => (x"c1",x"f0",x"ff",x"c0"),
   266 => (x"cd",x"f4",x"49",x"d1"),
   267 => (x"70",x"86",x"c4",x"87"),
   268 => (x"87",x"d2",x"05",x"98"),
   269 => (x"cc",x"1e",x"c0",x"c8"),
   270 => (x"e6",x"fd",x"49",x"66"),
   271 => (x"70",x"86",x"c4",x"87"),
   272 => (x"48",x"d0",x"ff",x"4b"),
   273 => (x"48",x"73",x"78",x"c2"),
   274 => (x"0e",x"87",x"eb",x"f3"),
   275 => (x"5d",x"5c",x"5b",x"5e"),
   276 => (x"c0",x"1e",x"c0",x"0e"),
   277 => (x"c9",x"c1",x"f0",x"ff"),
   278 => (x"87",x"de",x"f3",x"49"),
   279 => (x"df",x"c2",x"1e",x"d2"),
   280 => (x"fe",x"fc",x"49",x"d4"),
   281 => (x"c0",x"86",x"c8",x"87"),
   282 => (x"d2",x"84",x"c1",x"4c"),
   283 => (x"f8",x"04",x"ac",x"b7"),
   284 => (x"d4",x"df",x"c2",x"87"),
   285 => (x"c3",x"49",x"bf",x"97"),
   286 => (x"c0",x"c1",x"99",x"c0"),
   287 => (x"e7",x"c0",x"05",x"a9"),
   288 => (x"db",x"df",x"c2",x"87"),
   289 => (x"d0",x"49",x"bf",x"97"),
   290 => (x"dc",x"df",x"c2",x"31"),
   291 => (x"c8",x"4a",x"bf",x"97"),
   292 => (x"c2",x"b1",x"72",x"32"),
   293 => (x"bf",x"97",x"dd",x"df"),
   294 => (x"4c",x"71",x"b1",x"4a"),
   295 => (x"ff",x"ff",x"ff",x"cf"),
   296 => (x"ca",x"84",x"c1",x"9c"),
   297 => (x"87",x"e7",x"c1",x"34"),
   298 => (x"97",x"dd",x"df",x"c2"),
   299 => (x"31",x"c1",x"49",x"bf"),
   300 => (x"df",x"c2",x"99",x"c6"),
   301 => (x"4a",x"bf",x"97",x"de"),
   302 => (x"72",x"2a",x"b7",x"c7"),
   303 => (x"d9",x"df",x"c2",x"b1"),
   304 => (x"4d",x"4a",x"bf",x"97"),
   305 => (x"df",x"c2",x"9d",x"cf"),
   306 => (x"4a",x"bf",x"97",x"da"),
   307 => (x"32",x"ca",x"9a",x"c3"),
   308 => (x"97",x"db",x"df",x"c2"),
   309 => (x"33",x"c2",x"4b",x"bf"),
   310 => (x"df",x"c2",x"b2",x"73"),
   311 => (x"4b",x"bf",x"97",x"dc"),
   312 => (x"c6",x"9b",x"c0",x"c3"),
   313 => (x"b2",x"73",x"2b",x"b7"),
   314 => (x"48",x"c1",x"81",x"c2"),
   315 => (x"49",x"70",x"30",x"71"),
   316 => (x"30",x"75",x"48",x"c1"),
   317 => (x"4c",x"72",x"4d",x"70"),
   318 => (x"94",x"71",x"84",x"c1"),
   319 => (x"ad",x"b7",x"c0",x"c8"),
   320 => (x"c1",x"87",x"cc",x"06"),
   321 => (x"c8",x"2d",x"b7",x"34"),
   322 => (x"01",x"ad",x"b7",x"c0"),
   323 => (x"74",x"87",x"f4",x"ff"),
   324 => (x"87",x"de",x"f0",x"48"),
   325 => (x"5c",x"5b",x"5e",x"0e"),
   326 => (x"86",x"f8",x"0e",x"5d"),
   327 => (x"48",x"fa",x"e7",x"c2"),
   328 => (x"df",x"c2",x"78",x"c0"),
   329 => (x"49",x"c0",x"1e",x"f2"),
   330 => (x"c4",x"87",x"de",x"fb"),
   331 => (x"05",x"98",x"70",x"86"),
   332 => (x"48",x"c0",x"87",x"c5"),
   333 => (x"c0",x"87",x"ce",x"c9"),
   334 => (x"c0",x"7e",x"c1",x"4d"),
   335 => (x"49",x"bf",x"f6",x"f2"),
   336 => (x"4a",x"e8",x"e0",x"c2"),
   337 => (x"ec",x"4b",x"c8",x"71"),
   338 => (x"98",x"70",x"87",x"e0"),
   339 => (x"c0",x"87",x"c2",x"05"),
   340 => (x"f2",x"f2",x"c0",x"7e"),
   341 => (x"e1",x"c2",x"49",x"bf"),
   342 => (x"c8",x"71",x"4a",x"c4"),
   343 => (x"87",x"ca",x"ec",x"4b"),
   344 => (x"c2",x"05",x"98",x"70"),
   345 => (x"6e",x"7e",x"c0",x"87"),
   346 => (x"87",x"fd",x"c0",x"02"),
   347 => (x"bf",x"f8",x"e6",x"c2"),
   348 => (x"f0",x"e7",x"c2",x"4d"),
   349 => (x"48",x"7e",x"bf",x"9f"),
   350 => (x"a8",x"ea",x"d6",x"c5"),
   351 => (x"c2",x"87",x"c7",x"05"),
   352 => (x"4d",x"bf",x"f8",x"e6"),
   353 => (x"48",x"6e",x"87",x"ce"),
   354 => (x"a8",x"d5",x"e9",x"ca"),
   355 => (x"c0",x"87",x"c5",x"02"),
   356 => (x"87",x"f1",x"c7",x"48"),
   357 => (x"1e",x"f2",x"df",x"c2"),
   358 => (x"ec",x"f9",x"49",x"75"),
   359 => (x"70",x"86",x"c4",x"87"),
   360 => (x"87",x"c5",x"05",x"98"),
   361 => (x"dc",x"c7",x"48",x"c0"),
   362 => (x"f2",x"f2",x"c0",x"87"),
   363 => (x"e1",x"c2",x"49",x"bf"),
   364 => (x"c8",x"71",x"4a",x"c4"),
   365 => (x"87",x"f2",x"ea",x"4b"),
   366 => (x"c8",x"05",x"98",x"70"),
   367 => (x"fa",x"e7",x"c2",x"87"),
   368 => (x"da",x"78",x"c1",x"48"),
   369 => (x"f6",x"f2",x"c0",x"87"),
   370 => (x"e0",x"c2",x"49",x"bf"),
   371 => (x"c8",x"71",x"4a",x"e8"),
   372 => (x"87",x"d6",x"ea",x"4b"),
   373 => (x"c0",x"02",x"98",x"70"),
   374 => (x"48",x"c0",x"87",x"c5"),
   375 => (x"c2",x"87",x"e6",x"c6"),
   376 => (x"bf",x"97",x"f0",x"e7"),
   377 => (x"a9",x"d5",x"c1",x"49"),
   378 => (x"87",x"cd",x"c0",x"05"),
   379 => (x"97",x"f1",x"e7",x"c2"),
   380 => (x"ea",x"c2",x"49",x"bf"),
   381 => (x"c5",x"c0",x"02",x"a9"),
   382 => (x"c6",x"48",x"c0",x"87"),
   383 => (x"df",x"c2",x"87",x"c7"),
   384 => (x"7e",x"bf",x"97",x"f2"),
   385 => (x"a8",x"e9",x"c3",x"48"),
   386 => (x"87",x"ce",x"c0",x"02"),
   387 => (x"eb",x"c3",x"48",x"6e"),
   388 => (x"c5",x"c0",x"02",x"a8"),
   389 => (x"c5",x"48",x"c0",x"87"),
   390 => (x"df",x"c2",x"87",x"eb"),
   391 => (x"49",x"bf",x"97",x"fd"),
   392 => (x"cc",x"c0",x"05",x"99"),
   393 => (x"fe",x"df",x"c2",x"87"),
   394 => (x"c2",x"49",x"bf",x"97"),
   395 => (x"c5",x"c0",x"02",x"a9"),
   396 => (x"c5",x"48",x"c0",x"87"),
   397 => (x"df",x"c2",x"87",x"cf"),
   398 => (x"48",x"bf",x"97",x"ff"),
   399 => (x"58",x"f6",x"e7",x"c2"),
   400 => (x"c1",x"48",x"4c",x"70"),
   401 => (x"fa",x"e7",x"c2",x"88"),
   402 => (x"c0",x"e0",x"c2",x"58"),
   403 => (x"75",x"49",x"bf",x"97"),
   404 => (x"c1",x"e0",x"c2",x"81"),
   405 => (x"c8",x"4a",x"bf",x"97"),
   406 => (x"7e",x"a1",x"72",x"32"),
   407 => (x"48",x"c7",x"ec",x"c2"),
   408 => (x"e0",x"c2",x"78",x"6e"),
   409 => (x"48",x"bf",x"97",x"c2"),
   410 => (x"c2",x"58",x"a6",x"c8"),
   411 => (x"02",x"bf",x"fa",x"e7"),
   412 => (x"c0",x"87",x"d4",x"c2"),
   413 => (x"49",x"bf",x"f2",x"f2"),
   414 => (x"4a",x"c4",x"e1",x"c2"),
   415 => (x"e7",x"4b",x"c8",x"71"),
   416 => (x"98",x"70",x"87",x"e8"),
   417 => (x"87",x"c5",x"c0",x"02"),
   418 => (x"f8",x"c3",x"48",x"c0"),
   419 => (x"f2",x"e7",x"c2",x"87"),
   420 => (x"ec",x"c2",x"4c",x"bf"),
   421 => (x"e0",x"c2",x"5c",x"db"),
   422 => (x"49",x"bf",x"97",x"d7"),
   423 => (x"e0",x"c2",x"31",x"c8"),
   424 => (x"4a",x"bf",x"97",x"d6"),
   425 => (x"e0",x"c2",x"49",x"a1"),
   426 => (x"4a",x"bf",x"97",x"d8"),
   427 => (x"a1",x"72",x"32",x"d0"),
   428 => (x"d9",x"e0",x"c2",x"49"),
   429 => (x"d8",x"4a",x"bf",x"97"),
   430 => (x"49",x"a1",x"72",x"32"),
   431 => (x"c2",x"91",x"66",x"c4"),
   432 => (x"81",x"bf",x"c7",x"ec"),
   433 => (x"59",x"cf",x"ec",x"c2"),
   434 => (x"97",x"df",x"e0",x"c2"),
   435 => (x"32",x"c8",x"4a",x"bf"),
   436 => (x"97",x"de",x"e0",x"c2"),
   437 => (x"4a",x"a2",x"4b",x"bf"),
   438 => (x"97",x"e0",x"e0",x"c2"),
   439 => (x"33",x"d0",x"4b",x"bf"),
   440 => (x"c2",x"4a",x"a2",x"73"),
   441 => (x"bf",x"97",x"e1",x"e0"),
   442 => (x"d8",x"9b",x"cf",x"4b"),
   443 => (x"4a",x"a2",x"73",x"33"),
   444 => (x"5a",x"d3",x"ec",x"c2"),
   445 => (x"bf",x"cf",x"ec",x"c2"),
   446 => (x"74",x"8a",x"c2",x"4a"),
   447 => (x"d3",x"ec",x"c2",x"92"),
   448 => (x"78",x"a1",x"72",x"48"),
   449 => (x"c2",x"87",x"ca",x"c1"),
   450 => (x"bf",x"97",x"c4",x"e0"),
   451 => (x"c2",x"31",x"c8",x"49"),
   452 => (x"bf",x"97",x"c3",x"e0"),
   453 => (x"c2",x"49",x"a1",x"4a"),
   454 => (x"c2",x"59",x"c2",x"e8"),
   455 => (x"49",x"bf",x"fe",x"e7"),
   456 => (x"ff",x"c7",x"31",x"c5"),
   457 => (x"c2",x"29",x"c9",x"81"),
   458 => (x"c2",x"59",x"db",x"ec"),
   459 => (x"bf",x"97",x"c9",x"e0"),
   460 => (x"c2",x"32",x"c8",x"4a"),
   461 => (x"bf",x"97",x"c8",x"e0"),
   462 => (x"c4",x"4a",x"a2",x"4b"),
   463 => (x"82",x"6e",x"92",x"66"),
   464 => (x"5a",x"d7",x"ec",x"c2"),
   465 => (x"48",x"cf",x"ec",x"c2"),
   466 => (x"ec",x"c2",x"78",x"c0"),
   467 => (x"a1",x"72",x"48",x"cb"),
   468 => (x"db",x"ec",x"c2",x"78"),
   469 => (x"cf",x"ec",x"c2",x"48"),
   470 => (x"ec",x"c2",x"78",x"bf"),
   471 => (x"ec",x"c2",x"48",x"df"),
   472 => (x"c2",x"78",x"bf",x"d3"),
   473 => (x"02",x"bf",x"fa",x"e7"),
   474 => (x"74",x"87",x"c9",x"c0"),
   475 => (x"70",x"30",x"c4",x"48"),
   476 => (x"87",x"c9",x"c0",x"7e"),
   477 => (x"bf",x"d7",x"ec",x"c2"),
   478 => (x"70",x"30",x"c4",x"48"),
   479 => (x"fe",x"e7",x"c2",x"7e"),
   480 => (x"c1",x"78",x"6e",x"48"),
   481 => (x"26",x"8e",x"f8",x"48"),
   482 => (x"26",x"4c",x"26",x"4d"),
   483 => (x"0e",x"4f",x"26",x"4b"),
   484 => (x"5d",x"5c",x"5b",x"5e"),
   485 => (x"c2",x"4a",x"71",x"0e"),
   486 => (x"02",x"bf",x"fa",x"e7"),
   487 => (x"4b",x"72",x"87",x"cb"),
   488 => (x"4c",x"72",x"2b",x"c7"),
   489 => (x"c9",x"9c",x"ff",x"c1"),
   490 => (x"c8",x"4b",x"72",x"87"),
   491 => (x"c3",x"4c",x"72",x"2b"),
   492 => (x"ec",x"c2",x"9c",x"ff"),
   493 => (x"c0",x"83",x"bf",x"c7"),
   494 => (x"ab",x"bf",x"ee",x"f2"),
   495 => (x"c0",x"87",x"d9",x"02"),
   496 => (x"c2",x"5b",x"f2",x"f2"),
   497 => (x"73",x"1e",x"f2",x"df"),
   498 => (x"87",x"fd",x"f0",x"49"),
   499 => (x"98",x"70",x"86",x"c4"),
   500 => (x"c0",x"87",x"c5",x"05"),
   501 => (x"87",x"e6",x"c0",x"48"),
   502 => (x"bf",x"fa",x"e7",x"c2"),
   503 => (x"74",x"87",x"d2",x"02"),
   504 => (x"c2",x"91",x"c4",x"49"),
   505 => (x"69",x"81",x"f2",x"df"),
   506 => (x"ff",x"ff",x"cf",x"4d"),
   507 => (x"cb",x"9d",x"ff",x"ff"),
   508 => (x"c2",x"49",x"74",x"87"),
   509 => (x"f2",x"df",x"c2",x"91"),
   510 => (x"4d",x"69",x"9f",x"81"),
   511 => (x"c6",x"fe",x"48",x"75"),
   512 => (x"5b",x"5e",x"0e",x"87"),
   513 => (x"f8",x"0e",x"5d",x"5c"),
   514 => (x"9c",x"4c",x"71",x"86"),
   515 => (x"c0",x"87",x"c5",x"05"),
   516 => (x"87",x"c1",x"c3",x"48"),
   517 => (x"6e",x"7e",x"a4",x"c8"),
   518 => (x"d8",x"78",x"c0",x"48"),
   519 => (x"87",x"c7",x"02",x"66"),
   520 => (x"bf",x"97",x"66",x"d8"),
   521 => (x"c0",x"87",x"c5",x"05"),
   522 => (x"87",x"e9",x"c2",x"48"),
   523 => (x"49",x"c1",x"1e",x"c0"),
   524 => (x"c4",x"87",x"e0",x"ca"),
   525 => (x"9d",x"4d",x"70",x"86"),
   526 => (x"87",x"c2",x"c1",x"02"),
   527 => (x"4a",x"c2",x"e8",x"c2"),
   528 => (x"e0",x"49",x"66",x"d8"),
   529 => (x"98",x"70",x"87",x"c9"),
   530 => (x"87",x"f2",x"c0",x"02"),
   531 => (x"66",x"d8",x"4a",x"75"),
   532 => (x"e0",x"4b",x"cb",x"49"),
   533 => (x"98",x"70",x"87",x"ee"),
   534 => (x"87",x"e2",x"c0",x"02"),
   535 => (x"9d",x"75",x"1e",x"c0"),
   536 => (x"c8",x"87",x"c7",x"02"),
   537 => (x"78",x"c0",x"48",x"a6"),
   538 => (x"a6",x"c8",x"87",x"c5"),
   539 => (x"c8",x"78",x"c1",x"48"),
   540 => (x"de",x"c9",x"49",x"66"),
   541 => (x"70",x"86",x"c4",x"87"),
   542 => (x"fe",x"05",x"9d",x"4d"),
   543 => (x"9d",x"75",x"87",x"fe"),
   544 => (x"87",x"cf",x"c1",x"02"),
   545 => (x"6e",x"49",x"a5",x"dc"),
   546 => (x"da",x"78",x"69",x"48"),
   547 => (x"a6",x"c4",x"49",x"a5"),
   548 => (x"78",x"a4",x"c4",x"48"),
   549 => (x"c4",x"48",x"69",x"9f"),
   550 => (x"c2",x"78",x"08",x"66"),
   551 => (x"02",x"bf",x"fa",x"e7"),
   552 => (x"a5",x"d4",x"87",x"d2"),
   553 => (x"49",x"69",x"9f",x"49"),
   554 => (x"99",x"ff",x"ff",x"c0"),
   555 => (x"30",x"d0",x"48",x"71"),
   556 => (x"87",x"c2",x"7e",x"70"),
   557 => (x"49",x"6e",x"7e",x"c0"),
   558 => (x"bf",x"66",x"c4",x"48"),
   559 => (x"08",x"66",x"c4",x"80"),
   560 => (x"cc",x"7c",x"c0",x"78"),
   561 => (x"66",x"c4",x"49",x"a4"),
   562 => (x"a4",x"d0",x"79",x"bf"),
   563 => (x"c1",x"79",x"c0",x"49"),
   564 => (x"c0",x"87",x"c2",x"48"),
   565 => (x"fa",x"8e",x"f8",x"48"),
   566 => (x"5e",x"0e",x"87",x"ed"),
   567 => (x"0e",x"5d",x"5c",x"5b"),
   568 => (x"02",x"9c",x"4c",x"71"),
   569 => (x"c8",x"87",x"ca",x"c1"),
   570 => (x"02",x"69",x"49",x"a4"),
   571 => (x"d0",x"87",x"c2",x"c1"),
   572 => (x"49",x"6c",x"4a",x"66"),
   573 => (x"5a",x"a6",x"d4",x"82"),
   574 => (x"b9",x"4d",x"66",x"d0"),
   575 => (x"bf",x"f6",x"e7",x"c2"),
   576 => (x"72",x"ba",x"ff",x"4a"),
   577 => (x"02",x"99",x"71",x"99"),
   578 => (x"c4",x"87",x"e4",x"c0"),
   579 => (x"49",x"6b",x"4b",x"a4"),
   580 => (x"70",x"87",x"fc",x"f9"),
   581 => (x"f2",x"e7",x"c2",x"7b"),
   582 => (x"81",x"6c",x"49",x"bf"),
   583 => (x"b9",x"75",x"7c",x"71"),
   584 => (x"bf",x"f6",x"e7",x"c2"),
   585 => (x"72",x"ba",x"ff",x"4a"),
   586 => (x"05",x"99",x"71",x"99"),
   587 => (x"75",x"87",x"dc",x"ff"),
   588 => (x"87",x"d3",x"f9",x"7c"),
   589 => (x"71",x"1e",x"73",x"1e"),
   590 => (x"c7",x"02",x"9b",x"4b"),
   591 => (x"49",x"a3",x"c8",x"87"),
   592 => (x"87",x"c5",x"05",x"69"),
   593 => (x"f7",x"c0",x"48",x"c0"),
   594 => (x"cb",x"ec",x"c2",x"87"),
   595 => (x"a3",x"c4",x"4a",x"bf"),
   596 => (x"c2",x"49",x"69",x"49"),
   597 => (x"f2",x"e7",x"c2",x"89"),
   598 => (x"a2",x"71",x"91",x"bf"),
   599 => (x"f6",x"e7",x"c2",x"4a"),
   600 => (x"99",x"6b",x"49",x"bf"),
   601 => (x"c0",x"4a",x"a2",x"71"),
   602 => (x"c8",x"5a",x"f2",x"f2"),
   603 => (x"49",x"72",x"1e",x"66"),
   604 => (x"c4",x"87",x"d6",x"ea"),
   605 => (x"05",x"98",x"70",x"86"),
   606 => (x"48",x"c0",x"87",x"c4"),
   607 => (x"48",x"c1",x"87",x"c2"),
   608 => (x"1e",x"87",x"c8",x"f8"),
   609 => (x"4b",x"71",x"1e",x"73"),
   610 => (x"87",x"c7",x"02",x"9b"),
   611 => (x"69",x"49",x"a3",x"c8"),
   612 => (x"c0",x"87",x"c5",x"05"),
   613 => (x"87",x"f7",x"c0",x"48"),
   614 => (x"bf",x"cb",x"ec",x"c2"),
   615 => (x"49",x"a3",x"c4",x"4a"),
   616 => (x"89",x"c2",x"49",x"69"),
   617 => (x"bf",x"f2",x"e7",x"c2"),
   618 => (x"4a",x"a2",x"71",x"91"),
   619 => (x"bf",x"f6",x"e7",x"c2"),
   620 => (x"71",x"99",x"6b",x"49"),
   621 => (x"f2",x"c0",x"4a",x"a2"),
   622 => (x"66",x"c8",x"5a",x"f2"),
   623 => (x"e5",x"49",x"72",x"1e"),
   624 => (x"86",x"c4",x"87",x"ff"),
   625 => (x"c4",x"05",x"98",x"70"),
   626 => (x"c2",x"48",x"c0",x"87"),
   627 => (x"f6",x"48",x"c1",x"87"),
   628 => (x"5e",x"0e",x"87",x"f9"),
   629 => (x"1e",x"0e",x"5c",x"5b"),
   630 => (x"66",x"d0",x"4b",x"71"),
   631 => (x"73",x"2c",x"c9",x"4c"),
   632 => (x"d4",x"c1",x"02",x"9b"),
   633 => (x"49",x"a3",x"c8",x"87"),
   634 => (x"cc",x"c1",x"02",x"69"),
   635 => (x"f6",x"e7",x"c2",x"87"),
   636 => (x"b9",x"ff",x"49",x"bf"),
   637 => (x"7e",x"99",x"4a",x"6b"),
   638 => (x"d1",x"03",x"ac",x"71"),
   639 => (x"d0",x"7b",x"c0",x"87"),
   640 => (x"79",x"c0",x"49",x"a3"),
   641 => (x"c4",x"4a",x"a3",x"cc"),
   642 => (x"79",x"6a",x"49",x"a3"),
   643 => (x"8c",x"72",x"87",x"c2"),
   644 => (x"c0",x"02",x"9c",x"74"),
   645 => (x"1e",x"49",x"87",x"e3"),
   646 => (x"fd",x"fa",x"49",x"73"),
   647 => (x"d0",x"86",x"c4",x"87"),
   648 => (x"ff",x"c7",x"49",x"66"),
   649 => (x"87",x"cb",x"02",x"99"),
   650 => (x"1e",x"f2",x"df",x"c2"),
   651 => (x"c3",x"fc",x"49",x"73"),
   652 => (x"d0",x"86",x"c4",x"87"),
   653 => (x"66",x"d0",x"49",x"a3"),
   654 => (x"cc",x"f5",x"26",x"79"),
   655 => (x"1e",x"73",x"1e",x"87"),
   656 => (x"02",x"9b",x"4b",x"71"),
   657 => (x"c2",x"87",x"e4",x"c0"),
   658 => (x"73",x"5b",x"df",x"ec"),
   659 => (x"c2",x"8a",x"c2",x"4a"),
   660 => (x"49",x"bf",x"f2",x"e7"),
   661 => (x"cb",x"ec",x"c2",x"92"),
   662 => (x"80",x"72",x"48",x"bf"),
   663 => (x"58",x"e3",x"ec",x"c2"),
   664 => (x"30",x"c4",x"48",x"71"),
   665 => (x"58",x"c2",x"e8",x"c2"),
   666 => (x"c2",x"87",x"ed",x"c0"),
   667 => (x"c2",x"48",x"db",x"ec"),
   668 => (x"78",x"bf",x"cf",x"ec"),
   669 => (x"48",x"df",x"ec",x"c2"),
   670 => (x"bf",x"d3",x"ec",x"c2"),
   671 => (x"fa",x"e7",x"c2",x"78"),
   672 => (x"87",x"c9",x"02",x"bf"),
   673 => (x"bf",x"f2",x"e7",x"c2"),
   674 => (x"c7",x"31",x"c4",x"49"),
   675 => (x"d7",x"ec",x"c2",x"87"),
   676 => (x"31",x"c4",x"49",x"bf"),
   677 => (x"59",x"c2",x"e8",x"c2"),
   678 => (x"0e",x"87",x"f0",x"f3"),
   679 => (x"0e",x"5c",x"5b",x"5e"),
   680 => (x"4b",x"c0",x"4a",x"71"),
   681 => (x"c0",x"02",x"9a",x"72"),
   682 => (x"a2",x"da",x"87",x"e1"),
   683 => (x"4b",x"69",x"9f",x"49"),
   684 => (x"bf",x"fa",x"e7",x"c2"),
   685 => (x"d4",x"87",x"cf",x"02"),
   686 => (x"69",x"9f",x"49",x"a2"),
   687 => (x"ff",x"c0",x"4c",x"49"),
   688 => (x"34",x"d0",x"9c",x"ff"),
   689 => (x"4c",x"c0",x"87",x"c2"),
   690 => (x"73",x"b3",x"49",x"74"),
   691 => (x"87",x"ed",x"fd",x"49"),
   692 => (x"0e",x"87",x"f6",x"f2"),
   693 => (x"5d",x"5c",x"5b",x"5e"),
   694 => (x"71",x"86",x"f4",x"0e"),
   695 => (x"72",x"7e",x"c0",x"4a"),
   696 => (x"87",x"d8",x"02",x"9a"),
   697 => (x"48",x"ee",x"df",x"c2"),
   698 => (x"df",x"c2",x"78",x"c0"),
   699 => (x"ec",x"c2",x"48",x"e6"),
   700 => (x"c2",x"78",x"bf",x"df"),
   701 => (x"c2",x"48",x"ea",x"df"),
   702 => (x"78",x"bf",x"db",x"ec"),
   703 => (x"48",x"cf",x"e8",x"c2"),
   704 => (x"e7",x"c2",x"50",x"c0"),
   705 => (x"c2",x"49",x"bf",x"fe"),
   706 => (x"4a",x"bf",x"ee",x"df"),
   707 => (x"c4",x"03",x"aa",x"71"),
   708 => (x"49",x"72",x"87",x"c9"),
   709 => (x"c0",x"05",x"99",x"cf"),
   710 => (x"f2",x"c0",x"87",x"e9"),
   711 => (x"df",x"c2",x"48",x"ee"),
   712 => (x"c2",x"78",x"bf",x"e6"),
   713 => (x"c2",x"1e",x"f2",x"df"),
   714 => (x"49",x"bf",x"e6",x"df"),
   715 => (x"48",x"e6",x"df",x"c2"),
   716 => (x"71",x"78",x"a1",x"c1"),
   717 => (x"c4",x"87",x"d2",x"e3"),
   718 => (x"ea",x"f2",x"c0",x"86"),
   719 => (x"f2",x"df",x"c2",x"48"),
   720 => (x"c0",x"87",x"cc",x"78"),
   721 => (x"48",x"bf",x"ea",x"f2"),
   722 => (x"c0",x"80",x"e0",x"c0"),
   723 => (x"c2",x"58",x"ee",x"f2"),
   724 => (x"48",x"bf",x"ee",x"df"),
   725 => (x"df",x"c2",x"80",x"c1"),
   726 => (x"aa",x"27",x"58",x"f2"),
   727 => (x"bf",x"00",x"00",x"0c"),
   728 => (x"9d",x"4d",x"bf",x"97"),
   729 => (x"87",x"e3",x"c2",x"02"),
   730 => (x"02",x"ad",x"e5",x"c3"),
   731 => (x"c0",x"87",x"dc",x"c2"),
   732 => (x"4b",x"bf",x"ea",x"f2"),
   733 => (x"11",x"49",x"a3",x"cb"),
   734 => (x"05",x"ac",x"cf",x"4c"),
   735 => (x"75",x"87",x"d2",x"c1"),
   736 => (x"c1",x"99",x"df",x"49"),
   737 => (x"c2",x"91",x"cd",x"89"),
   738 => (x"c1",x"81",x"c2",x"e8"),
   739 => (x"51",x"12",x"4a",x"a3"),
   740 => (x"12",x"4a",x"a3",x"c3"),
   741 => (x"4a",x"a3",x"c5",x"51"),
   742 => (x"a3",x"c7",x"51",x"12"),
   743 => (x"c9",x"51",x"12",x"4a"),
   744 => (x"51",x"12",x"4a",x"a3"),
   745 => (x"12",x"4a",x"a3",x"ce"),
   746 => (x"4a",x"a3",x"d0",x"51"),
   747 => (x"a3",x"d2",x"51",x"12"),
   748 => (x"d4",x"51",x"12",x"4a"),
   749 => (x"51",x"12",x"4a",x"a3"),
   750 => (x"12",x"4a",x"a3",x"d6"),
   751 => (x"4a",x"a3",x"d8",x"51"),
   752 => (x"a3",x"dc",x"51",x"12"),
   753 => (x"de",x"51",x"12",x"4a"),
   754 => (x"51",x"12",x"4a",x"a3"),
   755 => (x"fa",x"c0",x"7e",x"c1"),
   756 => (x"c8",x"49",x"74",x"87"),
   757 => (x"eb",x"c0",x"05",x"99"),
   758 => (x"d0",x"49",x"74",x"87"),
   759 => (x"87",x"d1",x"05",x"99"),
   760 => (x"c0",x"02",x"66",x"dc"),
   761 => (x"49",x"73",x"87",x"cb"),
   762 => (x"70",x"0f",x"66",x"dc"),
   763 => (x"d3",x"c0",x"02",x"98"),
   764 => (x"c0",x"05",x"6e",x"87"),
   765 => (x"e8",x"c2",x"87",x"c6"),
   766 => (x"50",x"c0",x"48",x"c2"),
   767 => (x"bf",x"ea",x"f2",x"c0"),
   768 => (x"87",x"e1",x"c2",x"48"),
   769 => (x"48",x"cf",x"e8",x"c2"),
   770 => (x"c2",x"7e",x"50",x"c0"),
   771 => (x"49",x"bf",x"fe",x"e7"),
   772 => (x"bf",x"ee",x"df",x"c2"),
   773 => (x"04",x"aa",x"71",x"4a"),
   774 => (x"c2",x"87",x"f7",x"fb"),
   775 => (x"05",x"bf",x"df",x"ec"),
   776 => (x"c2",x"87",x"c8",x"c0"),
   777 => (x"02",x"bf",x"fa",x"e7"),
   778 => (x"c2",x"87",x"f8",x"c1"),
   779 => (x"49",x"bf",x"ea",x"df"),
   780 => (x"70",x"87",x"dc",x"ed"),
   781 => (x"ee",x"df",x"c2",x"49"),
   782 => (x"48",x"a6",x"c4",x"59"),
   783 => (x"bf",x"ea",x"df",x"c2"),
   784 => (x"fa",x"e7",x"c2",x"78"),
   785 => (x"d8",x"c0",x"02",x"bf"),
   786 => (x"49",x"66",x"c4",x"87"),
   787 => (x"ff",x"ff",x"ff",x"cf"),
   788 => (x"02",x"a9",x"99",x"f8"),
   789 => (x"c0",x"87",x"c5",x"c0"),
   790 => (x"87",x"e1",x"c0",x"4c"),
   791 => (x"dc",x"c0",x"4c",x"c1"),
   792 => (x"49",x"66",x"c4",x"87"),
   793 => (x"99",x"f8",x"ff",x"cf"),
   794 => (x"c8",x"c0",x"02",x"a9"),
   795 => (x"48",x"a6",x"c8",x"87"),
   796 => (x"c5",x"c0",x"78",x"c0"),
   797 => (x"48",x"a6",x"c8",x"87"),
   798 => (x"66",x"c8",x"78",x"c1"),
   799 => (x"05",x"9c",x"74",x"4c"),
   800 => (x"c4",x"87",x"e0",x"c0"),
   801 => (x"89",x"c2",x"49",x"66"),
   802 => (x"bf",x"f2",x"e7",x"c2"),
   803 => (x"ec",x"c2",x"91",x"4a"),
   804 => (x"c2",x"4a",x"bf",x"cb"),
   805 => (x"72",x"48",x"e6",x"df"),
   806 => (x"df",x"c2",x"78",x"a1"),
   807 => (x"78",x"c0",x"48",x"ee"),
   808 => (x"c0",x"87",x"df",x"f9"),
   809 => (x"eb",x"8e",x"f4",x"48"),
   810 => (x"00",x"00",x"87",x"dd"),
   811 => (x"ff",x"ff",x"00",x"00"),
   812 => (x"0c",x"ba",x"ff",x"ff"),
   813 => (x"0c",x"c3",x"00",x"00"),
   814 => (x"41",x"46",x"00",x"00"),
   815 => (x"20",x"32",x"33",x"54"),
   816 => (x"46",x"00",x"20",x"20"),
   817 => (x"36",x"31",x"54",x"41"),
   818 => (x"00",x"20",x"20",x"20"),
   819 => (x"48",x"d4",x"ff",x"1e"),
   820 => (x"68",x"78",x"ff",x"c3"),
   821 => (x"1e",x"4f",x"26",x"48"),
   822 => (x"c3",x"48",x"d4",x"ff"),
   823 => (x"d0",x"ff",x"78",x"ff"),
   824 => (x"78",x"e1",x"c0",x"48"),
   825 => (x"d4",x"48",x"d4",x"ff"),
   826 => (x"e3",x"ec",x"c2",x"78"),
   827 => (x"bf",x"d4",x"ff",x"48"),
   828 => (x"1e",x"4f",x"26",x"50"),
   829 => (x"c0",x"48",x"d0",x"ff"),
   830 => (x"4f",x"26",x"78",x"e0"),
   831 => (x"87",x"cc",x"ff",x"1e"),
   832 => (x"02",x"99",x"49",x"70"),
   833 => (x"fb",x"c0",x"87",x"c6"),
   834 => (x"87",x"f1",x"05",x"a9"),
   835 => (x"4f",x"26",x"48",x"71"),
   836 => (x"5c",x"5b",x"5e",x"0e"),
   837 => (x"c0",x"4b",x"71",x"0e"),
   838 => (x"87",x"f0",x"fe",x"4c"),
   839 => (x"02",x"99",x"49",x"70"),
   840 => (x"c0",x"87",x"f9",x"c0"),
   841 => (x"c0",x"02",x"a9",x"ec"),
   842 => (x"fb",x"c0",x"87",x"f2"),
   843 => (x"eb",x"c0",x"02",x"a9"),
   844 => (x"b7",x"66",x"cc",x"87"),
   845 => (x"87",x"c7",x"03",x"ac"),
   846 => (x"c2",x"02",x"66",x"d0"),
   847 => (x"71",x"53",x"71",x"87"),
   848 => (x"87",x"c2",x"02",x"99"),
   849 => (x"c3",x"fe",x"84",x"c1"),
   850 => (x"99",x"49",x"70",x"87"),
   851 => (x"c0",x"87",x"cd",x"02"),
   852 => (x"c7",x"02",x"a9",x"ec"),
   853 => (x"a9",x"fb",x"c0",x"87"),
   854 => (x"87",x"d5",x"ff",x"05"),
   855 => (x"c3",x"02",x"66",x"d0"),
   856 => (x"7b",x"97",x"c0",x"87"),
   857 => (x"05",x"a9",x"ec",x"c0"),
   858 => (x"4a",x"74",x"87",x"c4"),
   859 => (x"4a",x"74",x"87",x"c5"),
   860 => (x"72",x"8a",x"0a",x"c0"),
   861 => (x"26",x"87",x"c2",x"48"),
   862 => (x"26",x"4c",x"26",x"4d"),
   863 => (x"1e",x"4f",x"26",x"4b"),
   864 => (x"70",x"87",x"c9",x"fd"),
   865 => (x"f0",x"c0",x"4a",x"49"),
   866 => (x"87",x"c9",x"04",x"aa"),
   867 => (x"01",x"aa",x"f9",x"c0"),
   868 => (x"f0",x"c0",x"87",x"c3"),
   869 => (x"aa",x"c1",x"c1",x"8a"),
   870 => (x"c1",x"87",x"c9",x"04"),
   871 => (x"c3",x"01",x"aa",x"da"),
   872 => (x"8a",x"f7",x"c0",x"87"),
   873 => (x"04",x"aa",x"e1",x"c1"),
   874 => (x"fa",x"c1",x"87",x"c9"),
   875 => (x"87",x"c3",x"01",x"aa"),
   876 => (x"72",x"8a",x"fd",x"c0"),
   877 => (x"0e",x"4f",x"26",x"48"),
   878 => (x"0e",x"5c",x"5b",x"5e"),
   879 => (x"d4",x"ff",x"4a",x"71"),
   880 => (x"c0",x"49",x"72",x"4c"),
   881 => (x"4b",x"70",x"87",x"e9"),
   882 => (x"87",x"c2",x"02",x"9b"),
   883 => (x"d0",x"ff",x"8b",x"c1"),
   884 => (x"c1",x"78",x"c5",x"48"),
   885 => (x"49",x"73",x"7c",x"d5"),
   886 => (x"e3",x"c1",x"31",x"c6"),
   887 => (x"4a",x"bf",x"97",x"fa"),
   888 => (x"70",x"b0",x"71",x"48"),
   889 => (x"48",x"d0",x"ff",x"7c"),
   890 => (x"48",x"73",x"78",x"c4"),
   891 => (x"0e",x"87",x"ca",x"fe"),
   892 => (x"5d",x"5c",x"5b",x"5e"),
   893 => (x"71",x"86",x"f8",x"0e"),
   894 => (x"fb",x"7e",x"c0",x"4c"),
   895 => (x"4b",x"c0",x"87",x"d9"),
   896 => (x"97",x"dc",x"fa",x"c0"),
   897 => (x"a9",x"c0",x"49",x"bf"),
   898 => (x"fb",x"87",x"cf",x"04"),
   899 => (x"83",x"c1",x"87",x"ee"),
   900 => (x"97",x"dc",x"fa",x"c0"),
   901 => (x"06",x"ab",x"49",x"bf"),
   902 => (x"fa",x"c0",x"87",x"f1"),
   903 => (x"02",x"bf",x"97",x"dc"),
   904 => (x"e7",x"fa",x"87",x"cf"),
   905 => (x"99",x"49",x"70",x"87"),
   906 => (x"c0",x"87",x"c6",x"02"),
   907 => (x"f1",x"05",x"a9",x"ec"),
   908 => (x"fa",x"4b",x"c0",x"87"),
   909 => (x"4d",x"70",x"87",x"d6"),
   910 => (x"c8",x"87",x"d1",x"fa"),
   911 => (x"cb",x"fa",x"58",x"a6"),
   912 => (x"c1",x"4a",x"70",x"87"),
   913 => (x"49",x"a4",x"c8",x"83"),
   914 => (x"ad",x"49",x"69",x"97"),
   915 => (x"c0",x"87",x"c7",x"02"),
   916 => (x"c0",x"05",x"ad",x"ff"),
   917 => (x"a4",x"c9",x"87",x"e7"),
   918 => (x"49",x"69",x"97",x"49"),
   919 => (x"02",x"a9",x"66",x"c4"),
   920 => (x"c0",x"48",x"87",x"c7"),
   921 => (x"d4",x"05",x"a8",x"ff"),
   922 => (x"49",x"a4",x"ca",x"87"),
   923 => (x"aa",x"49",x"69",x"97"),
   924 => (x"c0",x"87",x"c6",x"02"),
   925 => (x"c4",x"05",x"aa",x"ff"),
   926 => (x"d0",x"7e",x"c1",x"87"),
   927 => (x"ad",x"ec",x"c0",x"87"),
   928 => (x"c0",x"87",x"c6",x"02"),
   929 => (x"c4",x"05",x"ad",x"fb"),
   930 => (x"c1",x"4b",x"c0",x"87"),
   931 => (x"fe",x"02",x"6e",x"7e"),
   932 => (x"de",x"f9",x"87",x"e1"),
   933 => (x"f8",x"48",x"73",x"87"),
   934 => (x"87",x"db",x"fb",x"8e"),
   935 => (x"5b",x"5e",x"0e",x"00"),
   936 => (x"f8",x"0e",x"5d",x"5c"),
   937 => (x"ff",x"4d",x"71",x"86"),
   938 => (x"1e",x"75",x"4b",x"d4"),
   939 => (x"49",x"e8",x"ec",x"c2"),
   940 => (x"c4",x"87",x"ce",x"e5"),
   941 => (x"02",x"98",x"70",x"86"),
   942 => (x"c4",x"87",x"cc",x"c4"),
   943 => (x"e3",x"c1",x"48",x"a6"),
   944 => (x"75",x"78",x"bf",x"fc"),
   945 => (x"87",x"ef",x"fb",x"49"),
   946 => (x"c5",x"48",x"d0",x"ff"),
   947 => (x"7b",x"d6",x"c1",x"78"),
   948 => (x"a2",x"75",x"4a",x"c0"),
   949 => (x"c1",x"7b",x"11",x"49"),
   950 => (x"aa",x"b7",x"cb",x"82"),
   951 => (x"cc",x"87",x"f3",x"04"),
   952 => (x"7b",x"ff",x"c3",x"4a"),
   953 => (x"e0",x"c0",x"82",x"c1"),
   954 => (x"f4",x"04",x"aa",x"b7"),
   955 => (x"48",x"d0",x"ff",x"87"),
   956 => (x"ff",x"c3",x"78",x"c4"),
   957 => (x"c1",x"78",x"c5",x"7b"),
   958 => (x"7b",x"c1",x"7b",x"d3"),
   959 => (x"48",x"66",x"78",x"c4"),
   960 => (x"06",x"a8",x"b7",x"c0"),
   961 => (x"c2",x"87",x"f0",x"c2"),
   962 => (x"4c",x"bf",x"f0",x"ec"),
   963 => (x"74",x"48",x"66",x"c4"),
   964 => (x"58",x"a6",x"c8",x"88"),
   965 => (x"c1",x"02",x"9c",x"74"),
   966 => (x"df",x"c2",x"87",x"f9"),
   967 => (x"c0",x"c8",x"7e",x"f2"),
   968 => (x"b7",x"c0",x"8c",x"4d"),
   969 => (x"87",x"c6",x"03",x"ac"),
   970 => (x"4d",x"a4",x"c0",x"c8"),
   971 => (x"ec",x"c2",x"4c",x"c0"),
   972 => (x"49",x"bf",x"97",x"e3"),
   973 => (x"d1",x"02",x"99",x"d0"),
   974 => (x"c2",x"1e",x"c0",x"87"),
   975 => (x"e7",x"49",x"e8",x"ec"),
   976 => (x"86",x"c4",x"87",x"f2"),
   977 => (x"c0",x"4a",x"49",x"70"),
   978 => (x"df",x"c2",x"87",x"ee"),
   979 => (x"ec",x"c2",x"1e",x"f2"),
   980 => (x"df",x"e7",x"49",x"e8"),
   981 => (x"70",x"86",x"c4",x"87"),
   982 => (x"d0",x"ff",x"4a",x"49"),
   983 => (x"78",x"c5",x"c8",x"48"),
   984 => (x"6e",x"7b",x"d4",x"c1"),
   985 => (x"6e",x"7b",x"bf",x"97"),
   986 => (x"70",x"80",x"c1",x"48"),
   987 => (x"05",x"8d",x"c1",x"7e"),
   988 => (x"ff",x"87",x"f0",x"ff"),
   989 => (x"78",x"c4",x"48",x"d0"),
   990 => (x"c5",x"05",x"9a",x"72"),
   991 => (x"c1",x"48",x"c0",x"87"),
   992 => (x"1e",x"c1",x"87",x"c7"),
   993 => (x"49",x"e8",x"ec",x"c2"),
   994 => (x"c4",x"87",x"cf",x"e5"),
   995 => (x"05",x"9c",x"74",x"86"),
   996 => (x"c4",x"87",x"c7",x"fe"),
   997 => (x"b7",x"c0",x"48",x"66"),
   998 => (x"87",x"d1",x"06",x"a8"),
   999 => (x"48",x"e8",x"ec",x"c2"),
  1000 => (x"80",x"d0",x"78",x"c0"),
  1001 => (x"80",x"f4",x"78",x"c0"),
  1002 => (x"bf",x"f4",x"ec",x"c2"),
  1003 => (x"48",x"66",x"c4",x"78"),
  1004 => (x"01",x"a8",x"b7",x"c0"),
  1005 => (x"ff",x"87",x"d0",x"fd"),
  1006 => (x"78",x"c5",x"48",x"d0"),
  1007 => (x"c0",x"7b",x"d3",x"c1"),
  1008 => (x"c1",x"78",x"c4",x"7b"),
  1009 => (x"c0",x"87",x"c2",x"48"),
  1010 => (x"26",x"8e",x"f8",x"48"),
  1011 => (x"26",x"4c",x"26",x"4d"),
  1012 => (x"0e",x"4f",x"26",x"4b"),
  1013 => (x"5d",x"5c",x"5b",x"5e"),
  1014 => (x"4b",x"71",x"1e",x"0e"),
  1015 => (x"ab",x"4d",x"4c",x"c0"),
  1016 => (x"87",x"e8",x"c0",x"04"),
  1017 => (x"1e",x"ef",x"f7",x"c0"),
  1018 => (x"c4",x"02",x"9d",x"75"),
  1019 => (x"c2",x"4a",x"c0",x"87"),
  1020 => (x"72",x"4a",x"c1",x"87"),
  1021 => (x"87",x"db",x"eb",x"49"),
  1022 => (x"7e",x"70",x"86",x"c4"),
  1023 => (x"05",x"6e",x"84",x"c1"),
  1024 => (x"4c",x"73",x"87",x"c2"),
  1025 => (x"ac",x"73",x"85",x"c1"),
  1026 => (x"87",x"d8",x"ff",x"06"),
  1027 => (x"fe",x"26",x"48",x"6e"),
  1028 => (x"5e",x"0e",x"87",x"f9"),
  1029 => (x"71",x"0e",x"5c",x"5b"),
  1030 => (x"02",x"66",x"cc",x"4b"),
  1031 => (x"c0",x"4c",x"87",x"d8"),
  1032 => (x"d8",x"02",x"8c",x"f0"),
  1033 => (x"c1",x"4a",x"74",x"87"),
  1034 => (x"87",x"d1",x"02",x"8a"),
  1035 => (x"87",x"cd",x"02",x"8a"),
  1036 => (x"87",x"c9",x"02",x"8a"),
  1037 => (x"49",x"73",x"87",x"d9"),
  1038 => (x"d2",x"87",x"e2",x"f9"),
  1039 => (x"c0",x"1e",x"74",x"87"),
  1040 => (x"d9",x"db",x"c1",x"49"),
  1041 => (x"73",x"1e",x"74",x"87"),
  1042 => (x"d1",x"db",x"c1",x"49"),
  1043 => (x"fd",x"86",x"c8",x"87"),
  1044 => (x"5e",x"0e",x"87",x"fb"),
  1045 => (x"0e",x"5d",x"5c",x"5b"),
  1046 => (x"49",x"4c",x"71",x"1e"),
  1047 => (x"ed",x"c2",x"91",x"de"),
  1048 => (x"85",x"71",x"4d",x"d0"),
  1049 => (x"c1",x"02",x"6d",x"97"),
  1050 => (x"ec",x"c2",x"87",x"dc"),
  1051 => (x"74",x"4a",x"bf",x"fc"),
  1052 => (x"fd",x"49",x"72",x"82"),
  1053 => (x"7e",x"70",x"87",x"dd"),
  1054 => (x"f2",x"c0",x"02",x"6e"),
  1055 => (x"c4",x"ed",x"c2",x"87"),
  1056 => (x"cb",x"4a",x"6e",x"4b"),
  1057 => (x"df",x"c0",x"ff",x"49"),
  1058 => (x"cb",x"4b",x"74",x"87"),
  1059 => (x"ce",x"e4",x"c1",x"93"),
  1060 => (x"c1",x"83",x"c4",x"83"),
  1061 => (x"74",x"7b",x"ca",x"c3"),
  1062 => (x"d1",x"c5",x"c1",x"49"),
  1063 => (x"c1",x"7b",x"75",x"87"),
  1064 => (x"bf",x"97",x"fb",x"e3"),
  1065 => (x"ed",x"c2",x"1e",x"49"),
  1066 => (x"e5",x"fd",x"49",x"c4"),
  1067 => (x"74",x"86",x"c4",x"87"),
  1068 => (x"f9",x"c4",x"c1",x"49"),
  1069 => (x"c1",x"49",x"c0",x"87"),
  1070 => (x"c2",x"87",x"d8",x"c6"),
  1071 => (x"c0",x"48",x"e4",x"ec"),
  1072 => (x"dd",x"49",x"c1",x"78"),
  1073 => (x"fc",x"26",x"87",x"d9"),
  1074 => (x"6f",x"4c",x"87",x"c1"),
  1075 => (x"6e",x"69",x"64",x"61"),
  1076 => (x"2e",x"2e",x"2e",x"67"),
  1077 => (x"5b",x"5e",x"0e",x"00"),
  1078 => (x"4b",x"71",x"0e",x"5c"),
  1079 => (x"fc",x"ec",x"c2",x"4a"),
  1080 => (x"49",x"72",x"82",x"bf"),
  1081 => (x"70",x"87",x"ec",x"fb"),
  1082 => (x"c4",x"02",x"9c",x"4c"),
  1083 => (x"ea",x"e6",x"49",x"87"),
  1084 => (x"fc",x"ec",x"c2",x"87"),
  1085 => (x"c1",x"78",x"c0",x"48"),
  1086 => (x"87",x"e3",x"dc",x"49"),
  1087 => (x"0e",x"87",x"ce",x"fb"),
  1088 => (x"5d",x"5c",x"5b",x"5e"),
  1089 => (x"c2",x"86",x"f4",x"0e"),
  1090 => (x"c0",x"4d",x"f2",x"df"),
  1091 => (x"48",x"a6",x"c4",x"4c"),
  1092 => (x"ec",x"c2",x"78",x"c0"),
  1093 => (x"c0",x"49",x"bf",x"fc"),
  1094 => (x"c1",x"c1",x"06",x"a9"),
  1095 => (x"f2",x"df",x"c2",x"87"),
  1096 => (x"c0",x"02",x"98",x"48"),
  1097 => (x"f7",x"c0",x"87",x"f8"),
  1098 => (x"66",x"c8",x"1e",x"ef"),
  1099 => (x"c4",x"87",x"c7",x"02"),
  1100 => (x"78",x"c0",x"48",x"a6"),
  1101 => (x"a6",x"c4",x"87",x"c5"),
  1102 => (x"c4",x"78",x"c1",x"48"),
  1103 => (x"d2",x"e6",x"49",x"66"),
  1104 => (x"70",x"86",x"c4",x"87"),
  1105 => (x"c4",x"84",x"c1",x"4d"),
  1106 => (x"80",x"c1",x"48",x"66"),
  1107 => (x"c2",x"58",x"a6",x"c8"),
  1108 => (x"49",x"bf",x"fc",x"ec"),
  1109 => (x"87",x"c6",x"03",x"ac"),
  1110 => (x"ff",x"05",x"9d",x"75"),
  1111 => (x"4c",x"c0",x"87",x"c8"),
  1112 => (x"c3",x"02",x"9d",x"75"),
  1113 => (x"f7",x"c0",x"87",x"e0"),
  1114 => (x"66",x"c8",x"1e",x"ef"),
  1115 => (x"cc",x"87",x"c7",x"02"),
  1116 => (x"78",x"c0",x"48",x"a6"),
  1117 => (x"a6",x"cc",x"87",x"c5"),
  1118 => (x"cc",x"78",x"c1",x"48"),
  1119 => (x"d2",x"e5",x"49",x"66"),
  1120 => (x"70",x"86",x"c4",x"87"),
  1121 => (x"c2",x"02",x"6e",x"7e"),
  1122 => (x"49",x"6e",x"87",x"e9"),
  1123 => (x"69",x"97",x"81",x"cb"),
  1124 => (x"02",x"99",x"d0",x"49"),
  1125 => (x"c1",x"87",x"d6",x"c1"),
  1126 => (x"74",x"4a",x"d5",x"c3"),
  1127 => (x"c1",x"91",x"cb",x"49"),
  1128 => (x"72",x"81",x"ce",x"e4"),
  1129 => (x"c3",x"81",x"c8",x"79"),
  1130 => (x"49",x"74",x"51",x"ff"),
  1131 => (x"ed",x"c2",x"91",x"de"),
  1132 => (x"85",x"71",x"4d",x"d0"),
  1133 => (x"7d",x"97",x"c1",x"c2"),
  1134 => (x"c0",x"49",x"a5",x"c1"),
  1135 => (x"e8",x"c2",x"51",x"e0"),
  1136 => (x"02",x"bf",x"97",x"c2"),
  1137 => (x"84",x"c1",x"87",x"d2"),
  1138 => (x"c2",x"4b",x"a5",x"c2"),
  1139 => (x"db",x"4a",x"c2",x"e8"),
  1140 => (x"d3",x"fb",x"fe",x"49"),
  1141 => (x"87",x"db",x"c1",x"87"),
  1142 => (x"c0",x"49",x"a5",x"cd"),
  1143 => (x"c2",x"84",x"c1",x"51"),
  1144 => (x"4a",x"6e",x"4b",x"a5"),
  1145 => (x"fa",x"fe",x"49",x"cb"),
  1146 => (x"c6",x"c1",x"87",x"fe"),
  1147 => (x"d2",x"c1",x"c1",x"87"),
  1148 => (x"cb",x"49",x"74",x"4a"),
  1149 => (x"ce",x"e4",x"c1",x"91"),
  1150 => (x"c2",x"79",x"72",x"81"),
  1151 => (x"bf",x"97",x"c2",x"e8"),
  1152 => (x"74",x"87",x"d8",x"02"),
  1153 => (x"c1",x"91",x"de",x"49"),
  1154 => (x"d0",x"ed",x"c2",x"84"),
  1155 => (x"c2",x"83",x"71",x"4b"),
  1156 => (x"dd",x"4a",x"c2",x"e8"),
  1157 => (x"cf",x"fa",x"fe",x"49"),
  1158 => (x"74",x"87",x"d8",x"87"),
  1159 => (x"c2",x"93",x"de",x"4b"),
  1160 => (x"cb",x"83",x"d0",x"ed"),
  1161 => (x"51",x"c0",x"49",x"a3"),
  1162 => (x"6e",x"73",x"84",x"c1"),
  1163 => (x"fe",x"49",x"cb",x"4a"),
  1164 => (x"c4",x"87",x"f5",x"f9"),
  1165 => (x"80",x"c1",x"48",x"66"),
  1166 => (x"c7",x"58",x"a6",x"c8"),
  1167 => (x"c5",x"c0",x"03",x"ac"),
  1168 => (x"fc",x"05",x"6e",x"87"),
  1169 => (x"48",x"74",x"87",x"e0"),
  1170 => (x"fe",x"f5",x"8e",x"f4"),
  1171 => (x"1e",x"73",x"1e",x"87"),
  1172 => (x"cb",x"49",x"4b",x"71"),
  1173 => (x"ce",x"e4",x"c1",x"91"),
  1174 => (x"4a",x"a1",x"c8",x"81"),
  1175 => (x"48",x"fa",x"e3",x"c1"),
  1176 => (x"a1",x"c9",x"50",x"12"),
  1177 => (x"dc",x"fa",x"c0",x"4a"),
  1178 => (x"ca",x"50",x"12",x"48"),
  1179 => (x"fb",x"e3",x"c1",x"81"),
  1180 => (x"c1",x"50",x"11",x"48"),
  1181 => (x"bf",x"97",x"fb",x"e3"),
  1182 => (x"49",x"c0",x"1e",x"49"),
  1183 => (x"c2",x"87",x"d3",x"f6"),
  1184 => (x"de",x"48",x"e4",x"ec"),
  1185 => (x"d6",x"49",x"c1",x"78"),
  1186 => (x"f5",x"26",x"87",x"d5"),
  1187 => (x"71",x"1e",x"87",x"c1"),
  1188 => (x"91",x"cb",x"49",x"4a"),
  1189 => (x"81",x"ce",x"e4",x"c1"),
  1190 => (x"48",x"11",x"81",x"c8"),
  1191 => (x"58",x"e8",x"ec",x"c2"),
  1192 => (x"48",x"fc",x"ec",x"c2"),
  1193 => (x"49",x"c1",x"78",x"c0"),
  1194 => (x"26",x"87",x"f4",x"d5"),
  1195 => (x"49",x"c0",x"1e",x"4f"),
  1196 => (x"87",x"df",x"fe",x"c0"),
  1197 => (x"71",x"1e",x"4f",x"26"),
  1198 => (x"87",x"d2",x"02",x"99"),
  1199 => (x"48",x"e3",x"e5",x"c1"),
  1200 => (x"80",x"f7",x"50",x"c0"),
  1201 => (x"40",x"ce",x"ca",x"c1"),
  1202 => (x"78",x"c7",x"e4",x"c1"),
  1203 => (x"e5",x"c1",x"87",x"ce"),
  1204 => (x"e4",x"c1",x"48",x"df"),
  1205 => (x"80",x"fc",x"78",x"c0"),
  1206 => (x"78",x"ed",x"ca",x"c1"),
  1207 => (x"5e",x"0e",x"4f",x"26"),
  1208 => (x"71",x"0e",x"5c",x"5b"),
  1209 => (x"92",x"cb",x"4a",x"4c"),
  1210 => (x"82",x"ce",x"e4",x"c1"),
  1211 => (x"c9",x"49",x"a2",x"c8"),
  1212 => (x"6b",x"97",x"4b",x"a2"),
  1213 => (x"69",x"97",x"1e",x"4b"),
  1214 => (x"82",x"ca",x"1e",x"49"),
  1215 => (x"e7",x"c0",x"49",x"12"),
  1216 => (x"49",x"c0",x"87",x"d8"),
  1217 => (x"74",x"87",x"d8",x"d4"),
  1218 => (x"e1",x"fb",x"c0",x"49"),
  1219 => (x"f2",x"8e",x"f8",x"87"),
  1220 => (x"73",x"1e",x"87",x"fb"),
  1221 => (x"49",x"4b",x"71",x"1e"),
  1222 => (x"73",x"87",x"c3",x"ff"),
  1223 => (x"87",x"fe",x"fe",x"49"),
  1224 => (x"1e",x"87",x"ec",x"f2"),
  1225 => (x"4b",x"71",x"1e",x"73"),
  1226 => (x"02",x"4a",x"a3",x"c6"),
  1227 => (x"8a",x"c1",x"87",x"db"),
  1228 => (x"8a",x"87",x"d6",x"02"),
  1229 => (x"87",x"da",x"c1",x"02"),
  1230 => (x"fc",x"c0",x"02",x"8a"),
  1231 => (x"c0",x"02",x"8a",x"87"),
  1232 => (x"02",x"8a",x"87",x"e1"),
  1233 => (x"db",x"c1",x"87",x"cb"),
  1234 => (x"fd",x"49",x"c7",x"87"),
  1235 => (x"de",x"c1",x"87",x"c0"),
  1236 => (x"fc",x"ec",x"c2",x"87"),
  1237 => (x"cb",x"c1",x"02",x"bf"),
  1238 => (x"88",x"c1",x"48",x"87"),
  1239 => (x"58",x"c0",x"ed",x"c2"),
  1240 => (x"c2",x"87",x"c1",x"c1"),
  1241 => (x"02",x"bf",x"c0",x"ed"),
  1242 => (x"c2",x"87",x"f9",x"c0"),
  1243 => (x"48",x"bf",x"fc",x"ec"),
  1244 => (x"ed",x"c2",x"80",x"c1"),
  1245 => (x"eb",x"c0",x"58",x"c0"),
  1246 => (x"fc",x"ec",x"c2",x"87"),
  1247 => (x"89",x"c6",x"49",x"bf"),
  1248 => (x"59",x"c0",x"ed",x"c2"),
  1249 => (x"03",x"a9",x"b7",x"c0"),
  1250 => (x"ec",x"c2",x"87",x"da"),
  1251 => (x"78",x"c0",x"48",x"fc"),
  1252 => (x"ed",x"c2",x"87",x"d2"),
  1253 => (x"cb",x"02",x"bf",x"c0"),
  1254 => (x"fc",x"ec",x"c2",x"87"),
  1255 => (x"80",x"c6",x"48",x"bf"),
  1256 => (x"58",x"c0",x"ed",x"c2"),
  1257 => (x"f6",x"d1",x"49",x"c0"),
  1258 => (x"c0",x"49",x"73",x"87"),
  1259 => (x"f0",x"87",x"ff",x"f8"),
  1260 => (x"5e",x"0e",x"87",x"dd"),
  1261 => (x"0e",x"5d",x"5c",x"5b"),
  1262 => (x"dc",x"86",x"d0",x"ff"),
  1263 => (x"a6",x"c8",x"59",x"a6"),
  1264 => (x"c4",x"78",x"c0",x"48"),
  1265 => (x"66",x"c4",x"c1",x"80"),
  1266 => (x"c1",x"80",x"c4",x"78"),
  1267 => (x"c1",x"80",x"c4",x"78"),
  1268 => (x"c0",x"ed",x"c2",x"78"),
  1269 => (x"c2",x"78",x"c1",x"48"),
  1270 => (x"48",x"bf",x"e4",x"ec"),
  1271 => (x"cb",x"05",x"a8",x"de"),
  1272 => (x"87",x"db",x"f4",x"87"),
  1273 => (x"a6",x"cc",x"49",x"70"),
  1274 => (x"87",x"f2",x"cf",x"59"),
  1275 => (x"e4",x"87",x"e8",x"e3"),
  1276 => (x"d7",x"e3",x"87",x"ca"),
  1277 => (x"c0",x"4c",x"70",x"87"),
  1278 => (x"c1",x"02",x"ac",x"fb"),
  1279 => (x"66",x"d8",x"87",x"fb"),
  1280 => (x"87",x"ed",x"c1",x"05"),
  1281 => (x"4a",x"66",x"c0",x"c1"),
  1282 => (x"7e",x"6a",x"82",x"c4"),
  1283 => (x"e0",x"c1",x"1e",x"72"),
  1284 => (x"66",x"c4",x"48",x"d3"),
  1285 => (x"4a",x"a1",x"c8",x"49"),
  1286 => (x"aa",x"71",x"41",x"20"),
  1287 => (x"10",x"87",x"f9",x"05"),
  1288 => (x"c1",x"4a",x"26",x"51"),
  1289 => (x"c1",x"48",x"66",x"c0"),
  1290 => (x"6a",x"78",x"cd",x"c9"),
  1291 => (x"74",x"81",x"c7",x"49"),
  1292 => (x"66",x"c0",x"c1",x"51"),
  1293 => (x"c1",x"81",x"c8",x"49"),
  1294 => (x"66",x"c0",x"c1",x"51"),
  1295 => (x"c0",x"81",x"c9",x"49"),
  1296 => (x"66",x"c0",x"c1",x"51"),
  1297 => (x"c0",x"81",x"ca",x"49"),
  1298 => (x"d8",x"1e",x"c1",x"51"),
  1299 => (x"c8",x"49",x"6a",x"1e"),
  1300 => (x"87",x"fc",x"e2",x"81"),
  1301 => (x"c4",x"c1",x"86",x"c8"),
  1302 => (x"a8",x"c0",x"48",x"66"),
  1303 => (x"c8",x"87",x"c7",x"01"),
  1304 => (x"78",x"c1",x"48",x"a6"),
  1305 => (x"c4",x"c1",x"87",x"ce"),
  1306 => (x"88",x"c1",x"48",x"66"),
  1307 => (x"c3",x"58",x"a6",x"d0"),
  1308 => (x"87",x"c8",x"e2",x"87"),
  1309 => (x"c2",x"48",x"a6",x"d0"),
  1310 => (x"02",x"9c",x"74",x"78"),
  1311 => (x"c8",x"87",x"db",x"cd"),
  1312 => (x"c8",x"c1",x"48",x"66"),
  1313 => (x"cd",x"03",x"a8",x"66"),
  1314 => (x"a6",x"dc",x"87",x"d0"),
  1315 => (x"e8",x"78",x"c0",x"48"),
  1316 => (x"e0",x"78",x"c0",x"80"),
  1317 => (x"4c",x"70",x"87",x"f6"),
  1318 => (x"05",x"ac",x"d0",x"c1"),
  1319 => (x"c4",x"87",x"d9",x"c2"),
  1320 => (x"da",x"e3",x"7e",x"66"),
  1321 => (x"c8",x"49",x"70",x"87"),
  1322 => (x"df",x"e0",x"59",x"a6"),
  1323 => (x"c0",x"4c",x"70",x"87"),
  1324 => (x"c1",x"05",x"ac",x"ec"),
  1325 => (x"66",x"c8",x"87",x"ed"),
  1326 => (x"c1",x"91",x"cb",x"49"),
  1327 => (x"c4",x"81",x"66",x"c0"),
  1328 => (x"4d",x"6a",x"4a",x"a1"),
  1329 => (x"c4",x"4a",x"a1",x"c8"),
  1330 => (x"ca",x"c1",x"52",x"66"),
  1331 => (x"df",x"ff",x"79",x"ce"),
  1332 => (x"4c",x"70",x"87",x"fa"),
  1333 => (x"87",x"d9",x"02",x"9c"),
  1334 => (x"02",x"ac",x"fb",x"c0"),
  1335 => (x"55",x"74",x"87",x"d3"),
  1336 => (x"87",x"e8",x"df",x"ff"),
  1337 => (x"02",x"9c",x"4c",x"70"),
  1338 => (x"fb",x"c0",x"87",x"c7"),
  1339 => (x"ed",x"ff",x"05",x"ac"),
  1340 => (x"55",x"e0",x"c0",x"87"),
  1341 => (x"c0",x"55",x"c1",x"c2"),
  1342 => (x"66",x"d8",x"7d",x"97"),
  1343 => (x"05",x"a9",x"6e",x"49"),
  1344 => (x"66",x"c8",x"87",x"db"),
  1345 => (x"a8",x"66",x"cc",x"48"),
  1346 => (x"c8",x"87",x"ca",x"04"),
  1347 => (x"80",x"c1",x"48",x"66"),
  1348 => (x"c8",x"58",x"a6",x"cc"),
  1349 => (x"48",x"66",x"cc",x"87"),
  1350 => (x"a6",x"d0",x"88",x"c1"),
  1351 => (x"eb",x"de",x"ff",x"58"),
  1352 => (x"c1",x"4c",x"70",x"87"),
  1353 => (x"c8",x"05",x"ac",x"d0"),
  1354 => (x"48",x"66",x"d4",x"87"),
  1355 => (x"a6",x"d8",x"80",x"c1"),
  1356 => (x"ac",x"d0",x"c1",x"58"),
  1357 => (x"87",x"e7",x"fd",x"02"),
  1358 => (x"48",x"a6",x"e0",x"c0"),
  1359 => (x"c4",x"78",x"66",x"d8"),
  1360 => (x"e0",x"c0",x"48",x"66"),
  1361 => (x"c9",x"05",x"a8",x"66"),
  1362 => (x"e4",x"c0",x"87",x"e2"),
  1363 => (x"78",x"c0",x"48",x"a6"),
  1364 => (x"78",x"c0",x"80",x"c4"),
  1365 => (x"fb",x"c0",x"48",x"74"),
  1366 => (x"6e",x"7e",x"70",x"88"),
  1367 => (x"87",x"e5",x"c8",x"02"),
  1368 => (x"88",x"cb",x"48",x"6e"),
  1369 => (x"02",x"6e",x"7e",x"70"),
  1370 => (x"6e",x"87",x"cd",x"c1"),
  1371 => (x"70",x"88",x"c9",x"48"),
  1372 => (x"c3",x"02",x"6e",x"7e"),
  1373 => (x"48",x"6e",x"87",x"e9"),
  1374 => (x"7e",x"70",x"88",x"c4"),
  1375 => (x"87",x"ce",x"02",x"6e"),
  1376 => (x"88",x"c1",x"48",x"6e"),
  1377 => (x"02",x"6e",x"7e",x"70"),
  1378 => (x"c7",x"87",x"d4",x"c3"),
  1379 => (x"a6",x"dc",x"87",x"f1"),
  1380 => (x"78",x"f0",x"c0",x"48"),
  1381 => (x"87",x"f4",x"dc",x"ff"),
  1382 => (x"ec",x"c0",x"4c",x"70"),
  1383 => (x"c4",x"c0",x"02",x"ac"),
  1384 => (x"a6",x"e0",x"c0",x"87"),
  1385 => (x"ac",x"ec",x"c0",x"5c"),
  1386 => (x"ff",x"87",x"cd",x"02"),
  1387 => (x"70",x"87",x"dd",x"dc"),
  1388 => (x"ac",x"ec",x"c0",x"4c"),
  1389 => (x"87",x"f3",x"ff",x"05"),
  1390 => (x"02",x"ac",x"ec",x"c0"),
  1391 => (x"ff",x"87",x"c4",x"c0"),
  1392 => (x"c0",x"87",x"c9",x"dc"),
  1393 => (x"d0",x"1e",x"ca",x"1e"),
  1394 => (x"91",x"cb",x"49",x"66"),
  1395 => (x"48",x"66",x"c8",x"c1"),
  1396 => (x"a6",x"cc",x"80",x"71"),
  1397 => (x"48",x"66",x"c8",x"58"),
  1398 => (x"a6",x"d0",x"80",x"c4"),
  1399 => (x"bf",x"66",x"cc",x"58"),
  1400 => (x"eb",x"dc",x"ff",x"49"),
  1401 => (x"de",x"1e",x"c1",x"87"),
  1402 => (x"bf",x"66",x"d4",x"1e"),
  1403 => (x"df",x"dc",x"ff",x"49"),
  1404 => (x"70",x"86",x"d0",x"87"),
  1405 => (x"89",x"09",x"c0",x"49"),
  1406 => (x"59",x"a6",x"ec",x"c0"),
  1407 => (x"48",x"66",x"e8",x"c0"),
  1408 => (x"c0",x"06",x"a8",x"c0"),
  1409 => (x"e8",x"c0",x"87",x"ee"),
  1410 => (x"a8",x"dd",x"48",x"66"),
  1411 => (x"87",x"e4",x"c0",x"03"),
  1412 => (x"49",x"bf",x"66",x"c4"),
  1413 => (x"81",x"66",x"e8",x"c0"),
  1414 => (x"c0",x"51",x"e0",x"c0"),
  1415 => (x"c1",x"49",x"66",x"e8"),
  1416 => (x"bf",x"66",x"c4",x"81"),
  1417 => (x"51",x"c1",x"c2",x"81"),
  1418 => (x"49",x"66",x"e8",x"c0"),
  1419 => (x"66",x"c4",x"81",x"c2"),
  1420 => (x"51",x"c0",x"81",x"bf"),
  1421 => (x"c9",x"c1",x"48",x"6e"),
  1422 => (x"49",x"6e",x"78",x"cd"),
  1423 => (x"66",x"d0",x"81",x"c8"),
  1424 => (x"c9",x"49",x"6e",x"51"),
  1425 => (x"51",x"66",x"d4",x"81"),
  1426 => (x"81",x"ca",x"49",x"6e"),
  1427 => (x"d0",x"51",x"66",x"dc"),
  1428 => (x"80",x"c1",x"48",x"66"),
  1429 => (x"48",x"58",x"a6",x"d4"),
  1430 => (x"78",x"c1",x"80",x"d8"),
  1431 => (x"ff",x"87",x"e6",x"c4"),
  1432 => (x"70",x"87",x"dc",x"dc"),
  1433 => (x"a6",x"ec",x"c0",x"49"),
  1434 => (x"d2",x"dc",x"ff",x"59"),
  1435 => (x"c0",x"49",x"70",x"87"),
  1436 => (x"dc",x"59",x"a6",x"e0"),
  1437 => (x"ec",x"c0",x"48",x"66"),
  1438 => (x"ca",x"c0",x"05",x"a8"),
  1439 => (x"48",x"a6",x"dc",x"87"),
  1440 => (x"78",x"66",x"e8",x"c0"),
  1441 => (x"ff",x"87",x"c4",x"c0"),
  1442 => (x"c8",x"87",x"c1",x"d9"),
  1443 => (x"91",x"cb",x"49",x"66"),
  1444 => (x"48",x"66",x"c0",x"c1"),
  1445 => (x"7e",x"70",x"80",x"71"),
  1446 => (x"81",x"c8",x"49",x"6e"),
  1447 => (x"82",x"ca",x"4a",x"6e"),
  1448 => (x"52",x"66",x"e8",x"c0"),
  1449 => (x"c1",x"4a",x"66",x"dc"),
  1450 => (x"66",x"e8",x"c0",x"82"),
  1451 => (x"72",x"48",x"c1",x"8a"),
  1452 => (x"c1",x"4a",x"70",x"30"),
  1453 => (x"79",x"97",x"72",x"8a"),
  1454 => (x"1e",x"49",x"69",x"97"),
  1455 => (x"49",x"66",x"ec",x"c0"),
  1456 => (x"c4",x"87",x"d9",x"d7"),
  1457 => (x"a6",x"f0",x"c0",x"86"),
  1458 => (x"c4",x"49",x"6e",x"58"),
  1459 => (x"c0",x"4d",x"69",x"81"),
  1460 => (x"c4",x"48",x"66",x"e0"),
  1461 => (x"c0",x"02",x"a8",x"66"),
  1462 => (x"a6",x"c4",x"87",x"c8"),
  1463 => (x"c0",x"78",x"c0",x"48"),
  1464 => (x"a6",x"c4",x"87",x"c5"),
  1465 => (x"c4",x"78",x"c1",x"48"),
  1466 => (x"e0",x"c0",x"1e",x"66"),
  1467 => (x"ff",x"49",x"75",x"1e"),
  1468 => (x"c8",x"87",x"dd",x"d8"),
  1469 => (x"c0",x"4c",x"70",x"86"),
  1470 => (x"c1",x"06",x"ac",x"b7"),
  1471 => (x"85",x"74",x"87",x"d4"),
  1472 => (x"74",x"49",x"e0",x"c0"),
  1473 => (x"c1",x"4b",x"75",x"89"),
  1474 => (x"71",x"4a",x"dc",x"e0"),
  1475 => (x"87",x"d8",x"e6",x"fe"),
  1476 => (x"e4",x"c0",x"85",x"c2"),
  1477 => (x"80",x"c1",x"48",x"66"),
  1478 => (x"58",x"a6",x"e8",x"c0"),
  1479 => (x"49",x"66",x"ec",x"c0"),
  1480 => (x"a9",x"70",x"81",x"c1"),
  1481 => (x"87",x"c8",x"c0",x"02"),
  1482 => (x"c0",x"48",x"a6",x"c4"),
  1483 => (x"87",x"c5",x"c0",x"78"),
  1484 => (x"c1",x"48",x"a6",x"c4"),
  1485 => (x"1e",x"66",x"c4",x"78"),
  1486 => (x"c0",x"49",x"a4",x"c2"),
  1487 => (x"88",x"71",x"48",x"e0"),
  1488 => (x"75",x"1e",x"49",x"70"),
  1489 => (x"c7",x"d7",x"ff",x"49"),
  1490 => (x"c0",x"86",x"c8",x"87"),
  1491 => (x"ff",x"01",x"a8",x"b7"),
  1492 => (x"e4",x"c0",x"87",x"c0"),
  1493 => (x"d1",x"c0",x"02",x"66"),
  1494 => (x"c9",x"49",x"6e",x"87"),
  1495 => (x"66",x"e4",x"c0",x"81"),
  1496 => (x"c1",x"48",x"6e",x"51"),
  1497 => (x"c0",x"78",x"de",x"cb"),
  1498 => (x"49",x"6e",x"87",x"cc"),
  1499 => (x"51",x"c2",x"81",x"c9"),
  1500 => (x"cc",x"c1",x"48",x"6e"),
  1501 => (x"e8",x"c0",x"78",x"d2"),
  1502 => (x"78",x"c1",x"48",x"a6"),
  1503 => (x"ff",x"87",x"c6",x"c0"),
  1504 => (x"70",x"87",x"f9",x"d5"),
  1505 => (x"66",x"e8",x"c0",x"4c"),
  1506 => (x"87",x"f5",x"c0",x"02"),
  1507 => (x"cc",x"48",x"66",x"c8"),
  1508 => (x"c0",x"04",x"a8",x"66"),
  1509 => (x"66",x"c8",x"87",x"cb"),
  1510 => (x"cc",x"80",x"c1",x"48"),
  1511 => (x"e0",x"c0",x"58",x"a6"),
  1512 => (x"48",x"66",x"cc",x"87"),
  1513 => (x"a6",x"d0",x"88",x"c1"),
  1514 => (x"87",x"d5",x"c0",x"58"),
  1515 => (x"05",x"ac",x"c6",x"c1"),
  1516 => (x"d0",x"87",x"c8",x"c0"),
  1517 => (x"80",x"c1",x"48",x"66"),
  1518 => (x"ff",x"58",x"a6",x"d4"),
  1519 => (x"70",x"87",x"fd",x"d4"),
  1520 => (x"48",x"66",x"d4",x"4c"),
  1521 => (x"a6",x"d8",x"80",x"c1"),
  1522 => (x"02",x"9c",x"74",x"58"),
  1523 => (x"c8",x"87",x"cb",x"c0"),
  1524 => (x"c8",x"c1",x"48",x"66"),
  1525 => (x"f2",x"04",x"a8",x"66"),
  1526 => (x"d4",x"ff",x"87",x"f0"),
  1527 => (x"66",x"c8",x"87",x"d5"),
  1528 => (x"03",x"a8",x"c7",x"48"),
  1529 => (x"c2",x"87",x"e5",x"c0"),
  1530 => (x"c0",x"48",x"c0",x"ed"),
  1531 => (x"49",x"66",x"c8",x"78"),
  1532 => (x"c0",x"c1",x"91",x"cb"),
  1533 => (x"a1",x"c4",x"81",x"66"),
  1534 => (x"c0",x"4a",x"6a",x"4a"),
  1535 => (x"66",x"c8",x"79",x"52"),
  1536 => (x"cc",x"80",x"c1",x"48"),
  1537 => (x"a8",x"c7",x"58",x"a6"),
  1538 => (x"87",x"db",x"ff",x"04"),
  1539 => (x"ff",x"8e",x"d0",x"ff"),
  1540 => (x"4c",x"87",x"f8",x"de"),
  1541 => (x"20",x"64",x"61",x"6f"),
  1542 => (x"00",x"20",x"2e",x"2a"),
  1543 => (x"1e",x"00",x"20",x"3a"),
  1544 => (x"4b",x"71",x"1e",x"73"),
  1545 => (x"87",x"c6",x"02",x"9b"),
  1546 => (x"48",x"fc",x"ec",x"c2"),
  1547 => (x"1e",x"c7",x"78",x"c0"),
  1548 => (x"bf",x"fc",x"ec",x"c2"),
  1549 => (x"e4",x"c1",x"1e",x"49"),
  1550 => (x"ec",x"c2",x"1e",x"ce"),
  1551 => (x"ed",x"49",x"bf",x"e4"),
  1552 => (x"86",x"cc",x"87",x"f0"),
  1553 => (x"bf",x"e4",x"ec",x"c2"),
  1554 => (x"87",x"ea",x"e9",x"49"),
  1555 => (x"c8",x"02",x"9b",x"73"),
  1556 => (x"ce",x"e4",x"c1",x"87"),
  1557 => (x"e7",x"e7",x"c0",x"49"),
  1558 => (x"f2",x"dd",x"ff",x"87"),
  1559 => (x"e3",x"c1",x"1e",x"87"),
  1560 => (x"50",x"c0",x"48",x"fa"),
  1561 => (x"bf",x"f1",x"e5",x"c1"),
  1562 => (x"f0",x"d8",x"ff",x"49"),
  1563 => (x"26",x"48",x"c0",x"87"),
  1564 => (x"e3",x"c7",x"1e",x"4f"),
  1565 => (x"fe",x"49",x"c1",x"87"),
  1566 => (x"e9",x"fe",x"87",x"e5"),
  1567 => (x"98",x"70",x"87",x"d2"),
  1568 => (x"fe",x"87",x"cd",x"02"),
  1569 => (x"70",x"87",x"cd",x"f2"),
  1570 => (x"87",x"c4",x"02",x"98"),
  1571 => (x"87",x"c2",x"4a",x"c1"),
  1572 => (x"9a",x"72",x"4a",x"c0"),
  1573 => (x"c0",x"87",x"ce",x"05"),
  1574 => (x"c1",x"e3",x"c1",x"1e"),
  1575 => (x"f7",x"f2",x"c0",x"49"),
  1576 => (x"fe",x"86",x"c4",x"87"),
  1577 => (x"c1",x"1e",x"c0",x"87"),
  1578 => (x"c0",x"49",x"cc",x"e3"),
  1579 => (x"c0",x"87",x"e9",x"f2"),
  1580 => (x"87",x"e9",x"fe",x"1e"),
  1581 => (x"f2",x"c0",x"49",x"70"),
  1582 => (x"da",x"c3",x"87",x"de"),
  1583 => (x"26",x"8e",x"f8",x"87"),
  1584 => (x"20",x"44",x"53",x"4f"),
  1585 => (x"6c",x"69",x"61",x"66"),
  1586 => (x"00",x"2e",x"64",x"65"),
  1587 => (x"74",x"6f",x"6f",x"42"),
  1588 => (x"2e",x"67",x"6e",x"69"),
  1589 => (x"1e",x"00",x"2e",x"2e"),
  1590 => (x"87",x"c0",x"ea",x"c0"),
  1591 => (x"87",x"ee",x"f5",x"c0"),
  1592 => (x"4f",x"26",x"87",x"f6"),
  1593 => (x"fc",x"ec",x"c2",x"1e"),
  1594 => (x"c2",x"78",x"c0",x"48"),
  1595 => (x"c0",x"48",x"e4",x"ec"),
  1596 => (x"87",x"fd",x"fd",x"78"),
  1597 => (x"48",x"c0",x"87",x"e1"),
  1598 => (x"00",x"00",x"4f",x"26"),
  1599 => (x"00",x"00",x"00",x"01"),
  1600 => (x"78",x"45",x"20",x"80"),
  1601 => (x"80",x"00",x"74",x"69"),
  1602 => (x"63",x"61",x"42",x"20"),
  1603 => (x"12",x"8e",x"00",x"6b"),
  1604 => (x"2b",x"50",x"00",x"00"),
  1605 => (x"00",x"00",x"00",x"00"),
  1606 => (x"00",x"12",x"8e",x"00"),
  1607 => (x"00",x"2b",x"6e",x"00"),
  1608 => (x"00",x"00",x"00",x"00"),
  1609 => (x"00",x"00",x"12",x"8e"),
  1610 => (x"00",x"00",x"2b",x"8c"),
  1611 => (x"8e",x"00",x"00",x"00"),
  1612 => (x"aa",x"00",x"00",x"12"),
  1613 => (x"00",x"00",x"00",x"2b"),
  1614 => (x"12",x"8e",x"00",x"00"),
  1615 => (x"2b",x"c8",x"00",x"00"),
  1616 => (x"00",x"00",x"00",x"00"),
  1617 => (x"00",x"12",x"8e",x"00"),
  1618 => (x"00",x"2b",x"e6",x"00"),
  1619 => (x"00",x"00",x"00",x"00"),
  1620 => (x"00",x"00",x"12",x"8e"),
  1621 => (x"00",x"00",x"2c",x"04"),
  1622 => (x"8e",x"00",x"00",x"00"),
  1623 => (x"00",x"00",x"00",x"12"),
  1624 => (x"00",x"00",x"00",x"00"),
  1625 => (x"13",x"23",x"00",x"00"),
  1626 => (x"00",x"00",x"00",x"00"),
  1627 => (x"00",x"00",x"00",x"00"),
  1628 => (x"00",x"19",x"75",x"00"),
  1629 => (x"34",x"36",x"43",x"00"),
  1630 => (x"20",x"20",x"20",x"20"),
  1631 => (x"4d",x"4f",x"52",x"20"),
  1632 => (x"f0",x"fe",x"1e",x"00"),
  1633 => (x"cd",x"78",x"c0",x"48"),
  1634 => (x"26",x"09",x"79",x"09"),
  1635 => (x"fe",x"1e",x"1e",x"4f"),
  1636 => (x"48",x"7e",x"bf",x"f0"),
  1637 => (x"1e",x"4f",x"26",x"26"),
  1638 => (x"c1",x"48",x"f0",x"fe"),
  1639 => (x"1e",x"4f",x"26",x"78"),
  1640 => (x"c0",x"48",x"f0",x"fe"),
  1641 => (x"1e",x"4f",x"26",x"78"),
  1642 => (x"52",x"c0",x"4a",x"71"),
  1643 => (x"0e",x"4f",x"26",x"52"),
  1644 => (x"5d",x"5c",x"5b",x"5e"),
  1645 => (x"71",x"86",x"f4",x"0e"),
  1646 => (x"7e",x"6d",x"97",x"4d"),
  1647 => (x"97",x"4c",x"a5",x"c1"),
  1648 => (x"a6",x"c8",x"48",x"6c"),
  1649 => (x"c4",x"48",x"6e",x"58"),
  1650 => (x"c5",x"05",x"a8",x"66"),
  1651 => (x"c0",x"48",x"ff",x"87"),
  1652 => (x"ca",x"ff",x"87",x"e6"),
  1653 => (x"49",x"a5",x"c2",x"87"),
  1654 => (x"71",x"4b",x"6c",x"97"),
  1655 => (x"6b",x"97",x"4b",x"a3"),
  1656 => (x"7e",x"6c",x"97",x"4b"),
  1657 => (x"80",x"c1",x"48",x"6e"),
  1658 => (x"c7",x"58",x"a6",x"c8"),
  1659 => (x"58",x"a6",x"cc",x"98"),
  1660 => (x"fe",x"7c",x"97",x"70"),
  1661 => (x"48",x"73",x"87",x"e1"),
  1662 => (x"4d",x"26",x"8e",x"f4"),
  1663 => (x"4b",x"26",x"4c",x"26"),
  1664 => (x"5e",x"0e",x"4f",x"26"),
  1665 => (x"f4",x"0e",x"5c",x"5b"),
  1666 => (x"d8",x"4c",x"71",x"86"),
  1667 => (x"ff",x"c3",x"4a",x"66"),
  1668 => (x"4b",x"a4",x"c2",x"9a"),
  1669 => (x"73",x"49",x"6c",x"97"),
  1670 => (x"51",x"72",x"49",x"a1"),
  1671 => (x"6e",x"7e",x"6c",x"97"),
  1672 => (x"c8",x"80",x"c1",x"48"),
  1673 => (x"98",x"c7",x"58",x"a6"),
  1674 => (x"70",x"58",x"a6",x"cc"),
  1675 => (x"ff",x"8e",x"f4",x"54"),
  1676 => (x"1e",x"1e",x"87",x"ca"),
  1677 => (x"e0",x"87",x"e8",x"fd"),
  1678 => (x"c0",x"49",x"4a",x"bf"),
  1679 => (x"02",x"99",x"c0",x"e0"),
  1680 => (x"1e",x"72",x"87",x"cb"),
  1681 => (x"49",x"e2",x"f0",x"c2"),
  1682 => (x"c4",x"87",x"f7",x"fe"),
  1683 => (x"87",x"fd",x"fc",x"86"),
  1684 => (x"c2",x"fd",x"7e",x"70"),
  1685 => (x"4f",x"26",x"26",x"87"),
  1686 => (x"e2",x"f0",x"c2",x"1e"),
  1687 => (x"87",x"c7",x"fd",x"49"),
  1688 => (x"49",x"f2",x"e8",x"c1"),
  1689 => (x"c4",x"87",x"da",x"fc"),
  1690 => (x"4f",x"26",x"87",x"c7"),
  1691 => (x"48",x"d0",x"ff",x"1e"),
  1692 => (x"ff",x"78",x"e1",x"c8"),
  1693 => (x"78",x"c5",x"48",x"d4"),
  1694 => (x"c3",x"02",x"66",x"c4"),
  1695 => (x"78",x"e0",x"c3",x"87"),
  1696 => (x"c6",x"02",x"66",x"c8"),
  1697 => (x"48",x"d4",x"ff",x"87"),
  1698 => (x"ff",x"78",x"f0",x"c3"),
  1699 => (x"78",x"71",x"48",x"d4"),
  1700 => (x"c8",x"48",x"d0",x"ff"),
  1701 => (x"e0",x"c0",x"78",x"e1"),
  1702 => (x"0e",x"4f",x"26",x"78"),
  1703 => (x"0e",x"5c",x"5b",x"5e"),
  1704 => (x"f0",x"c2",x"4c",x"71"),
  1705 => (x"c6",x"fc",x"49",x"e2"),
  1706 => (x"c0",x"4a",x"70",x"87"),
  1707 => (x"c2",x"04",x"aa",x"b7"),
  1708 => (x"f0",x"c3",x"87",x"e2"),
  1709 => (x"87",x"c9",x"05",x"aa"),
  1710 => (x"48",x"e0",x"ed",x"c1"),
  1711 => (x"c3",x"c2",x"78",x"c1"),
  1712 => (x"aa",x"e0",x"c3",x"87"),
  1713 => (x"c1",x"87",x"c9",x"05"),
  1714 => (x"c1",x"48",x"e4",x"ed"),
  1715 => (x"87",x"f4",x"c1",x"78"),
  1716 => (x"bf",x"e4",x"ed",x"c1"),
  1717 => (x"c2",x"87",x"c6",x"02"),
  1718 => (x"c2",x"4b",x"a2",x"c0"),
  1719 => (x"74",x"4b",x"72",x"87"),
  1720 => (x"87",x"d1",x"05",x"9c"),
  1721 => (x"bf",x"e0",x"ed",x"c1"),
  1722 => (x"e4",x"ed",x"c1",x"1e"),
  1723 => (x"49",x"72",x"1e",x"bf"),
  1724 => (x"c8",x"87",x"f9",x"fd"),
  1725 => (x"e0",x"ed",x"c1",x"86"),
  1726 => (x"e0",x"c0",x"02",x"bf"),
  1727 => (x"c4",x"49",x"73",x"87"),
  1728 => (x"c1",x"91",x"29",x"b7"),
  1729 => (x"73",x"81",x"c0",x"ef"),
  1730 => (x"c2",x"9a",x"cf",x"4a"),
  1731 => (x"72",x"48",x"c1",x"92"),
  1732 => (x"ff",x"4a",x"70",x"30"),
  1733 => (x"69",x"48",x"72",x"ba"),
  1734 => (x"db",x"79",x"70",x"98"),
  1735 => (x"c4",x"49",x"73",x"87"),
  1736 => (x"c1",x"91",x"29",x"b7"),
  1737 => (x"73",x"81",x"c0",x"ef"),
  1738 => (x"c2",x"9a",x"cf",x"4a"),
  1739 => (x"72",x"48",x"c3",x"92"),
  1740 => (x"48",x"4a",x"70",x"30"),
  1741 => (x"79",x"70",x"b0",x"69"),
  1742 => (x"48",x"e4",x"ed",x"c1"),
  1743 => (x"ed",x"c1",x"78",x"c0"),
  1744 => (x"78",x"c0",x"48",x"e0"),
  1745 => (x"49",x"e2",x"f0",x"c2"),
  1746 => (x"70",x"87",x"e4",x"f9"),
  1747 => (x"aa",x"b7",x"c0",x"4a"),
  1748 => (x"87",x"de",x"fd",x"03"),
  1749 => (x"87",x"c2",x"48",x"c0"),
  1750 => (x"4c",x"26",x"4d",x"26"),
  1751 => (x"4f",x"26",x"4b",x"26"),
  1752 => (x"00",x"00",x"00",x"00"),
  1753 => (x"00",x"00",x"00",x"00"),
  1754 => (x"49",x"4a",x"71",x"1e"),
  1755 => (x"26",x"87",x"ec",x"fc"),
  1756 => (x"4a",x"c0",x"1e",x"4f"),
  1757 => (x"91",x"c4",x"49",x"72"),
  1758 => (x"81",x"c0",x"ef",x"c1"),
  1759 => (x"82",x"c1",x"79",x"c0"),
  1760 => (x"04",x"aa",x"b7",x"d0"),
  1761 => (x"4f",x"26",x"87",x"ee"),
  1762 => (x"5c",x"5b",x"5e",x"0e"),
  1763 => (x"4d",x"71",x"0e",x"5d"),
  1764 => (x"75",x"87",x"cc",x"f8"),
  1765 => (x"2a",x"b7",x"c4",x"4a"),
  1766 => (x"c0",x"ef",x"c1",x"92"),
  1767 => (x"cf",x"4c",x"75",x"82"),
  1768 => (x"6a",x"94",x"c2",x"9c"),
  1769 => (x"2b",x"74",x"4b",x"49"),
  1770 => (x"48",x"c2",x"9b",x"c3"),
  1771 => (x"4c",x"70",x"30",x"74"),
  1772 => (x"48",x"74",x"bc",x"ff"),
  1773 => (x"7a",x"70",x"98",x"71"),
  1774 => (x"73",x"87",x"dc",x"f7"),
  1775 => (x"87",x"d8",x"fe",x"48"),
  1776 => (x"00",x"00",x"00",x"00"),
  1777 => (x"00",x"00",x"00",x"00"),
  1778 => (x"00",x"00",x"00",x"00"),
  1779 => (x"00",x"00",x"00",x"00"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"00",x"00",x"00",x"00"),
  1784 => (x"00",x"00",x"00",x"00"),
  1785 => (x"00",x"00",x"00",x"00"),
  1786 => (x"00",x"00",x"00",x"00"),
  1787 => (x"00",x"00",x"00",x"00"),
  1788 => (x"00",x"00",x"00",x"00"),
  1789 => (x"00",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"48",x"d0",x"ff",x"1e"),
  1793 => (x"71",x"78",x"e1",x"c8"),
  1794 => (x"08",x"d4",x"ff",x"48"),
  1795 => (x"1e",x"4f",x"26",x"78"),
  1796 => (x"c8",x"48",x"d0",x"ff"),
  1797 => (x"48",x"71",x"78",x"e1"),
  1798 => (x"78",x"08",x"d4",x"ff"),
  1799 => (x"ff",x"48",x"66",x"c4"),
  1800 => (x"26",x"78",x"08",x"d4"),
  1801 => (x"4a",x"71",x"1e",x"4f"),
  1802 => (x"1e",x"49",x"66",x"c4"),
  1803 => (x"de",x"ff",x"49",x"72"),
  1804 => (x"48",x"d0",x"ff",x"87"),
  1805 => (x"26",x"78",x"e0",x"c0"),
  1806 => (x"73",x"1e",x"4f",x"26"),
  1807 => (x"c8",x"4b",x"71",x"1e"),
  1808 => (x"73",x"1e",x"49",x"66"),
  1809 => (x"a2",x"e0",x"c1",x"4a"),
  1810 => (x"87",x"d9",x"ff",x"49"),
  1811 => (x"26",x"87",x"c4",x"26"),
  1812 => (x"26",x"4c",x"26",x"4d"),
  1813 => (x"1e",x"4f",x"26",x"4b"),
  1814 => (x"c3",x"4a",x"d4",x"ff"),
  1815 => (x"d0",x"ff",x"7a",x"ff"),
  1816 => (x"78",x"e1",x"c0",x"48"),
  1817 => (x"f0",x"c2",x"7a",x"de"),
  1818 => (x"49",x"7a",x"bf",x"ec"),
  1819 => (x"70",x"28",x"c8",x"48"),
  1820 => (x"d0",x"48",x"71",x"7a"),
  1821 => (x"71",x"7a",x"70",x"28"),
  1822 => (x"70",x"28",x"d8",x"48"),
  1823 => (x"f0",x"f0",x"c2",x"7a"),
  1824 => (x"48",x"49",x"7a",x"bf"),
  1825 => (x"7a",x"70",x"28",x"c8"),
  1826 => (x"28",x"d0",x"48",x"71"),
  1827 => (x"48",x"71",x"7a",x"70"),
  1828 => (x"7a",x"70",x"28",x"d8"),
  1829 => (x"c0",x"48",x"d0",x"ff"),
  1830 => (x"4f",x"26",x"78",x"e0"),
  1831 => (x"71",x"1e",x"73",x"1e"),
  1832 => (x"ec",x"f0",x"c2",x"4a"),
  1833 => (x"2b",x"72",x"4b",x"bf"),
  1834 => (x"04",x"aa",x"e0",x"c0"),
  1835 => (x"49",x"72",x"87",x"ce"),
  1836 => (x"c2",x"89",x"e0",x"c0"),
  1837 => (x"4b",x"bf",x"f0",x"f0"),
  1838 => (x"87",x"cf",x"2b",x"71"),
  1839 => (x"72",x"49",x"e0",x"c0"),
  1840 => (x"f0",x"f0",x"c2",x"89"),
  1841 => (x"30",x"71",x"48",x"bf"),
  1842 => (x"c8",x"b3",x"49",x"70"),
  1843 => (x"48",x"73",x"9b",x"66"),
  1844 => (x"4d",x"26",x"87",x"c4"),
  1845 => (x"4b",x"26",x"4c",x"26"),
  1846 => (x"5e",x"0e",x"4f",x"26"),
  1847 => (x"0e",x"5d",x"5c",x"5b"),
  1848 => (x"4b",x"71",x"86",x"ec"),
  1849 => (x"bf",x"ec",x"f0",x"c2"),
  1850 => (x"2c",x"73",x"4c",x"7e"),
  1851 => (x"04",x"ab",x"e0",x"c0"),
  1852 => (x"c4",x"87",x"e0",x"c0"),
  1853 => (x"78",x"c0",x"48",x"a6"),
  1854 => (x"e0",x"c0",x"49",x"73"),
  1855 => (x"c0",x"4a",x"71",x"89"),
  1856 => (x"72",x"48",x"66",x"e4"),
  1857 => (x"58",x"a6",x"cc",x"30"),
  1858 => (x"bf",x"f0",x"f0",x"c2"),
  1859 => (x"2c",x"71",x"4c",x"4d"),
  1860 => (x"73",x"87",x"e4",x"c0"),
  1861 => (x"66",x"e4",x"c0",x"49"),
  1862 => (x"c8",x"30",x"71",x"48"),
  1863 => (x"e0",x"c0",x"58",x"a6"),
  1864 => (x"c0",x"89",x"73",x"49"),
  1865 => (x"71",x"48",x"66",x"e4"),
  1866 => (x"58",x"a6",x"cc",x"28"),
  1867 => (x"bf",x"f0",x"f0",x"c2"),
  1868 => (x"30",x"71",x"48",x"4d"),
  1869 => (x"c0",x"b4",x"49",x"70"),
  1870 => (x"c1",x"9c",x"66",x"e4"),
  1871 => (x"66",x"e8",x"c0",x"84"),
  1872 => (x"87",x"c2",x"04",x"ac"),
  1873 => (x"e0",x"c0",x"4c",x"c0"),
  1874 => (x"87",x"d3",x"04",x"ab"),
  1875 => (x"c0",x"48",x"a6",x"cc"),
  1876 => (x"c0",x"49",x"73",x"78"),
  1877 => (x"48",x"74",x"89",x"e0"),
  1878 => (x"a6",x"d4",x"30",x"71"),
  1879 => (x"73",x"87",x"d5",x"58"),
  1880 => (x"71",x"48",x"74",x"49"),
  1881 => (x"58",x"a6",x"d0",x"30"),
  1882 => (x"73",x"49",x"e0",x"c0"),
  1883 => (x"71",x"48",x"74",x"89"),
  1884 => (x"58",x"a6",x"d4",x"28"),
  1885 => (x"ff",x"4a",x"66",x"c4"),
  1886 => (x"c8",x"9a",x"6e",x"ba"),
  1887 => (x"b9",x"ff",x"49",x"66"),
  1888 => (x"48",x"72",x"99",x"75"),
  1889 => (x"c2",x"b0",x"66",x"cc"),
  1890 => (x"71",x"58",x"f0",x"f0"),
  1891 => (x"b0",x"66",x"d0",x"48"),
  1892 => (x"58",x"f4",x"f0",x"c2"),
  1893 => (x"ec",x"87",x"c0",x"fb"),
  1894 => (x"87",x"f6",x"fc",x"8e"),
  1895 => (x"48",x"d0",x"ff",x"1e"),
  1896 => (x"71",x"78",x"c9",x"c8"),
  1897 => (x"08",x"d4",x"ff",x"48"),
  1898 => (x"1e",x"4f",x"26",x"78"),
  1899 => (x"eb",x"49",x"4a",x"71"),
  1900 => (x"48",x"d0",x"ff",x"87"),
  1901 => (x"4f",x"26",x"78",x"c8"),
  1902 => (x"71",x"1e",x"73",x"1e"),
  1903 => (x"c0",x"f1",x"c2",x"4b"),
  1904 => (x"87",x"c3",x"02",x"bf"),
  1905 => (x"ff",x"87",x"eb",x"c2"),
  1906 => (x"c9",x"c8",x"48",x"d0"),
  1907 => (x"c0",x"49",x"73",x"78"),
  1908 => (x"d4",x"ff",x"b1",x"e0"),
  1909 => (x"c2",x"78",x"71",x"48"),
  1910 => (x"c0",x"48",x"f4",x"f0"),
  1911 => (x"02",x"66",x"c8",x"78"),
  1912 => (x"ff",x"c3",x"87",x"c5"),
  1913 => (x"c0",x"87",x"c2",x"49"),
  1914 => (x"fc",x"f0",x"c2",x"49"),
  1915 => (x"02",x"66",x"cc",x"59"),
  1916 => (x"d5",x"c5",x"87",x"c6"),
  1917 => (x"87",x"c4",x"4a",x"d5"),
  1918 => (x"4a",x"ff",x"ff",x"cf"),
  1919 => (x"5a",x"c0",x"f1",x"c2"),
  1920 => (x"48",x"c0",x"f1",x"c2"),
  1921 => (x"87",x"c4",x"78",x"c1"),
  1922 => (x"4c",x"26",x"4d",x"26"),
  1923 => (x"4f",x"26",x"4b",x"26"),
  1924 => (x"5c",x"5b",x"5e",x"0e"),
  1925 => (x"4a",x"71",x"0e",x"5d"),
  1926 => (x"bf",x"fc",x"f0",x"c2"),
  1927 => (x"02",x"9a",x"72",x"4c"),
  1928 => (x"c8",x"49",x"87",x"cb"),
  1929 => (x"ee",x"f6",x"c1",x"91"),
  1930 => (x"c4",x"83",x"71",x"4b"),
  1931 => (x"ee",x"fa",x"c1",x"87"),
  1932 => (x"13",x"4d",x"c0",x"4b"),
  1933 => (x"c2",x"99",x"74",x"49"),
  1934 => (x"b9",x"bf",x"f8",x"f0"),
  1935 => (x"71",x"48",x"d4",x"ff"),
  1936 => (x"2c",x"b7",x"c1",x"78"),
  1937 => (x"ad",x"b7",x"c8",x"85"),
  1938 => (x"c2",x"87",x"e8",x"04"),
  1939 => (x"48",x"bf",x"f4",x"f0"),
  1940 => (x"f0",x"c2",x"80",x"c8"),
  1941 => (x"ef",x"fe",x"58",x"f8"),
  1942 => (x"1e",x"73",x"1e",x"87"),
  1943 => (x"4a",x"13",x"4b",x"71"),
  1944 => (x"87",x"cb",x"02",x"9a"),
  1945 => (x"e7",x"fe",x"49",x"72"),
  1946 => (x"9a",x"4a",x"13",x"87"),
  1947 => (x"fe",x"87",x"f5",x"05"),
  1948 => (x"c2",x"1e",x"87",x"da"),
  1949 => (x"49",x"bf",x"f4",x"f0"),
  1950 => (x"48",x"f4",x"f0",x"c2"),
  1951 => (x"c4",x"78",x"a1",x"c1"),
  1952 => (x"03",x"a9",x"b7",x"c0"),
  1953 => (x"d4",x"ff",x"87",x"db"),
  1954 => (x"f8",x"f0",x"c2",x"48"),
  1955 => (x"f0",x"c2",x"78",x"bf"),
  1956 => (x"c2",x"49",x"bf",x"f4"),
  1957 => (x"c1",x"48",x"f4",x"f0"),
  1958 => (x"c0",x"c4",x"78",x"a1"),
  1959 => (x"e5",x"04",x"a9",x"b7"),
  1960 => (x"48",x"d0",x"ff",x"87"),
  1961 => (x"f1",x"c2",x"78",x"c8"),
  1962 => (x"78",x"c0",x"48",x"c0"),
  1963 => (x"00",x"00",x"4f",x"26"),
  1964 => (x"00",x"00",x"00",x"00"),
  1965 => (x"00",x"00",x"00",x"00"),
  1966 => (x"00",x"5f",x"5f",x"00"),
  1967 => (x"03",x"00",x"00",x"00"),
  1968 => (x"03",x"03",x"00",x"03"),
  1969 => (x"7f",x"14",x"00",x"00"),
  1970 => (x"7f",x"7f",x"14",x"7f"),
  1971 => (x"24",x"00",x"00",x"14"),
  1972 => (x"3a",x"6b",x"6b",x"2e"),
  1973 => (x"6a",x"4c",x"00",x"12"),
  1974 => (x"56",x"6c",x"18",x"36"),
  1975 => (x"7e",x"30",x"00",x"32"),
  1976 => (x"3a",x"77",x"59",x"4f"),
  1977 => (x"00",x"00",x"40",x"68"),
  1978 => (x"00",x"03",x"07",x"04"),
  1979 => (x"00",x"00",x"00",x"00"),
  1980 => (x"41",x"63",x"3e",x"1c"),
  1981 => (x"00",x"00",x"00",x"00"),
  1982 => (x"1c",x"3e",x"63",x"41"),
  1983 => (x"2a",x"08",x"00",x"00"),
  1984 => (x"3e",x"1c",x"1c",x"3e"),
  1985 => (x"08",x"00",x"08",x"2a"),
  1986 => (x"08",x"3e",x"3e",x"08"),
  1987 => (x"00",x"00",x"00",x"08"),
  1988 => (x"00",x"60",x"e0",x"80"),
  1989 => (x"08",x"00",x"00",x"00"),
  1990 => (x"08",x"08",x"08",x"08"),
  1991 => (x"00",x"00",x"00",x"08"),
  1992 => (x"00",x"60",x"60",x"00"),
  1993 => (x"60",x"40",x"00",x"00"),
  1994 => (x"06",x"0c",x"18",x"30"),
  1995 => (x"3e",x"00",x"01",x"03"),
  1996 => (x"7f",x"4d",x"59",x"7f"),
  1997 => (x"04",x"00",x"00",x"3e"),
  1998 => (x"00",x"7f",x"7f",x"06"),
  1999 => (x"42",x"00",x"00",x"00"),
  2000 => (x"4f",x"59",x"71",x"63"),
  2001 => (x"22",x"00",x"00",x"46"),
  2002 => (x"7f",x"49",x"49",x"63"),
  2003 => (x"1c",x"18",x"00",x"36"),
  2004 => (x"7f",x"7f",x"13",x"16"),
  2005 => (x"27",x"00",x"00",x"10"),
  2006 => (x"7d",x"45",x"45",x"67"),
  2007 => (x"3c",x"00",x"00",x"39"),
  2008 => (x"79",x"49",x"4b",x"7e"),
  2009 => (x"01",x"00",x"00",x"30"),
  2010 => (x"0f",x"79",x"71",x"01"),
  2011 => (x"36",x"00",x"00",x"07"),
  2012 => (x"7f",x"49",x"49",x"7f"),
  2013 => (x"06",x"00",x"00",x"36"),
  2014 => (x"3f",x"69",x"49",x"4f"),
  2015 => (x"00",x"00",x"00",x"1e"),
  2016 => (x"00",x"66",x"66",x"00"),
  2017 => (x"00",x"00",x"00",x"00"),
  2018 => (x"00",x"66",x"e6",x"80"),
  2019 => (x"08",x"00",x"00",x"00"),
  2020 => (x"22",x"14",x"14",x"08"),
  2021 => (x"14",x"00",x"00",x"22"),
  2022 => (x"14",x"14",x"14",x"14"),
  2023 => (x"22",x"00",x"00",x"14"),
  2024 => (x"08",x"14",x"14",x"22"),
  2025 => (x"02",x"00",x"00",x"08"),
  2026 => (x"0f",x"59",x"51",x"03"),
  2027 => (x"7f",x"3e",x"00",x"06"),
  2028 => (x"1f",x"55",x"5d",x"41"),
  2029 => (x"7e",x"00",x"00",x"1e"),
  2030 => (x"7f",x"09",x"09",x"7f"),
  2031 => (x"7f",x"00",x"00",x"7e"),
  2032 => (x"7f",x"49",x"49",x"7f"),
  2033 => (x"1c",x"00",x"00",x"36"),
  2034 => (x"41",x"41",x"63",x"3e"),
  2035 => (x"7f",x"00",x"00",x"41"),
  2036 => (x"3e",x"63",x"41",x"7f"),
  2037 => (x"7f",x"00",x"00",x"1c"),
  2038 => (x"41",x"49",x"49",x"7f"),
  2039 => (x"7f",x"00",x"00",x"41"),
  2040 => (x"01",x"09",x"09",x"7f"),
  2041 => (x"3e",x"00",x"00",x"01"),
  2042 => (x"7b",x"49",x"41",x"7f"),
  2043 => (x"7f",x"00",x"00",x"7a"),
  2044 => (x"7f",x"08",x"08",x"7f"),
  2045 => (x"00",x"00",x"00",x"7f"),
  2046 => (x"41",x"7f",x"7f",x"41"),
  2047 => (x"20",x"00",x"00",x"00"),
  2048 => (x"7f",x"40",x"40",x"60"),
  2049 => (x"7f",x"7f",x"00",x"3f"),
  2050 => (x"63",x"36",x"1c",x"08"),
  2051 => (x"7f",x"00",x"00",x"41"),
  2052 => (x"40",x"40",x"40",x"7f"),
  2053 => (x"7f",x"7f",x"00",x"40"),
  2054 => (x"7f",x"06",x"0c",x"06"),
  2055 => (x"7f",x"7f",x"00",x"7f"),
  2056 => (x"7f",x"18",x"0c",x"06"),
  2057 => (x"3e",x"00",x"00",x"7f"),
  2058 => (x"7f",x"41",x"41",x"7f"),
  2059 => (x"7f",x"00",x"00",x"3e"),
  2060 => (x"0f",x"09",x"09",x"7f"),
  2061 => (x"7f",x"3e",x"00",x"06"),
  2062 => (x"7e",x"7f",x"61",x"41"),
  2063 => (x"7f",x"00",x"00",x"40"),
  2064 => (x"7f",x"19",x"09",x"7f"),
  2065 => (x"26",x"00",x"00",x"66"),
  2066 => (x"7b",x"59",x"4d",x"6f"),
  2067 => (x"01",x"00",x"00",x"32"),
  2068 => (x"01",x"7f",x"7f",x"01"),
  2069 => (x"3f",x"00",x"00",x"01"),
  2070 => (x"7f",x"40",x"40",x"7f"),
  2071 => (x"0f",x"00",x"00",x"3f"),
  2072 => (x"3f",x"70",x"70",x"3f"),
  2073 => (x"7f",x"7f",x"00",x"0f"),
  2074 => (x"7f",x"30",x"18",x"30"),
  2075 => (x"63",x"41",x"00",x"7f"),
  2076 => (x"36",x"1c",x"1c",x"36"),
  2077 => (x"03",x"01",x"41",x"63"),
  2078 => (x"06",x"7c",x"7c",x"06"),
  2079 => (x"71",x"61",x"01",x"03"),
  2080 => (x"43",x"47",x"4d",x"59"),
  2081 => (x"00",x"00",x"00",x"41"),
  2082 => (x"41",x"41",x"7f",x"7f"),
  2083 => (x"03",x"01",x"00",x"00"),
  2084 => (x"30",x"18",x"0c",x"06"),
  2085 => (x"00",x"00",x"40",x"60"),
  2086 => (x"7f",x"7f",x"41",x"41"),
  2087 => (x"0c",x"08",x"00",x"00"),
  2088 => (x"0c",x"06",x"03",x"06"),
  2089 => (x"80",x"80",x"00",x"08"),
  2090 => (x"80",x"80",x"80",x"80"),
  2091 => (x"00",x"00",x"00",x"80"),
  2092 => (x"04",x"07",x"03",x"00"),
  2093 => (x"20",x"00",x"00",x"00"),
  2094 => (x"7c",x"54",x"54",x"74"),
  2095 => (x"7f",x"00",x"00",x"78"),
  2096 => (x"7c",x"44",x"44",x"7f"),
  2097 => (x"38",x"00",x"00",x"38"),
  2098 => (x"44",x"44",x"44",x"7c"),
  2099 => (x"38",x"00",x"00",x"00"),
  2100 => (x"7f",x"44",x"44",x"7c"),
  2101 => (x"38",x"00",x"00",x"7f"),
  2102 => (x"5c",x"54",x"54",x"7c"),
  2103 => (x"04",x"00",x"00",x"18"),
  2104 => (x"05",x"05",x"7f",x"7e"),
  2105 => (x"18",x"00",x"00",x"00"),
  2106 => (x"fc",x"a4",x"a4",x"bc"),
  2107 => (x"7f",x"00",x"00",x"7c"),
  2108 => (x"7c",x"04",x"04",x"7f"),
  2109 => (x"00",x"00",x"00",x"78"),
  2110 => (x"40",x"7d",x"3d",x"00"),
  2111 => (x"80",x"00",x"00",x"00"),
  2112 => (x"7d",x"fd",x"80",x"80"),
  2113 => (x"7f",x"00",x"00",x"00"),
  2114 => (x"6c",x"38",x"10",x"7f"),
  2115 => (x"00",x"00",x"00",x"44"),
  2116 => (x"40",x"7f",x"3f",x"00"),
  2117 => (x"7c",x"7c",x"00",x"00"),
  2118 => (x"7c",x"0c",x"18",x"0c"),
  2119 => (x"7c",x"00",x"00",x"78"),
  2120 => (x"7c",x"04",x"04",x"7c"),
  2121 => (x"38",x"00",x"00",x"78"),
  2122 => (x"7c",x"44",x"44",x"7c"),
  2123 => (x"fc",x"00",x"00",x"38"),
  2124 => (x"3c",x"24",x"24",x"fc"),
  2125 => (x"18",x"00",x"00",x"18"),
  2126 => (x"fc",x"24",x"24",x"3c"),
  2127 => (x"7c",x"00",x"00",x"fc"),
  2128 => (x"0c",x"04",x"04",x"7c"),
  2129 => (x"48",x"00",x"00",x"08"),
  2130 => (x"74",x"54",x"54",x"5c"),
  2131 => (x"04",x"00",x"00",x"20"),
  2132 => (x"44",x"44",x"7f",x"3f"),
  2133 => (x"3c",x"00",x"00",x"00"),
  2134 => (x"7c",x"40",x"40",x"7c"),
  2135 => (x"1c",x"00",x"00",x"7c"),
  2136 => (x"3c",x"60",x"60",x"3c"),
  2137 => (x"7c",x"3c",x"00",x"1c"),
  2138 => (x"7c",x"60",x"30",x"60"),
  2139 => (x"6c",x"44",x"00",x"3c"),
  2140 => (x"6c",x"38",x"10",x"38"),
  2141 => (x"1c",x"00",x"00",x"44"),
  2142 => (x"3c",x"60",x"e0",x"bc"),
  2143 => (x"44",x"00",x"00",x"1c"),
  2144 => (x"4c",x"5c",x"74",x"64"),
  2145 => (x"08",x"00",x"00",x"44"),
  2146 => (x"41",x"77",x"3e",x"08"),
  2147 => (x"00",x"00",x"00",x"41"),
  2148 => (x"00",x"7f",x"7f",x"00"),
  2149 => (x"41",x"00",x"00",x"00"),
  2150 => (x"08",x"3e",x"77",x"41"),
  2151 => (x"01",x"02",x"00",x"08"),
  2152 => (x"02",x"02",x"03",x"01"),
  2153 => (x"7f",x"7f",x"00",x"01"),
  2154 => (x"7f",x"7f",x"7f",x"7f"),
  2155 => (x"08",x"08",x"00",x"7f"),
  2156 => (x"3e",x"3e",x"1c",x"1c"),
  2157 => (x"7f",x"7f",x"7f",x"7f"),
  2158 => (x"1c",x"1c",x"3e",x"3e"),
  2159 => (x"10",x"00",x"08",x"08"),
  2160 => (x"18",x"7c",x"7c",x"18"),
  2161 => (x"10",x"00",x"00",x"10"),
  2162 => (x"30",x"7c",x"7c",x"30"),
  2163 => (x"30",x"10",x"00",x"10"),
  2164 => (x"1e",x"78",x"60",x"60"),
  2165 => (x"66",x"42",x"00",x"06"),
  2166 => (x"66",x"3c",x"18",x"3c"),
  2167 => (x"38",x"78",x"00",x"42"),
  2168 => (x"6c",x"c6",x"c2",x"6a"),
  2169 => (x"00",x"60",x"00",x"38"),
  2170 => (x"00",x"00",x"60",x"00"),
  2171 => (x"5e",x"0e",x"00",x"60"),
  2172 => (x"0e",x"5d",x"5c",x"5b"),
  2173 => (x"c2",x"4c",x"71",x"1e"),
  2174 => (x"4d",x"bf",x"d1",x"f1"),
  2175 => (x"1e",x"c0",x"4b",x"c0"),
  2176 => (x"c7",x"02",x"ab",x"74"),
  2177 => (x"48",x"a6",x"c4",x"87"),
  2178 => (x"87",x"c5",x"78",x"c0"),
  2179 => (x"c1",x"48",x"a6",x"c4"),
  2180 => (x"1e",x"66",x"c4",x"78"),
  2181 => (x"df",x"ee",x"49",x"73"),
  2182 => (x"c0",x"86",x"c8",x"87"),
  2183 => (x"ef",x"ef",x"49",x"e0"),
  2184 => (x"4a",x"a5",x"c4",x"87"),
  2185 => (x"f0",x"f0",x"49",x"6a"),
  2186 => (x"87",x"c6",x"f1",x"87"),
  2187 => (x"83",x"c1",x"85",x"cb"),
  2188 => (x"04",x"ab",x"b7",x"c8"),
  2189 => (x"26",x"87",x"c7",x"ff"),
  2190 => (x"4c",x"26",x"4d",x"26"),
  2191 => (x"4f",x"26",x"4b",x"26"),
  2192 => (x"c2",x"4a",x"71",x"1e"),
  2193 => (x"c2",x"5a",x"d5",x"f1"),
  2194 => (x"c7",x"48",x"d5",x"f1"),
  2195 => (x"dd",x"fe",x"49",x"78"),
  2196 => (x"1e",x"4f",x"26",x"87"),
  2197 => (x"4a",x"71",x"1e",x"73"),
  2198 => (x"03",x"aa",x"b7",x"c0"),
  2199 => (x"d6",x"c2",x"87",x"d3"),
  2200 => (x"c4",x"05",x"bf",x"ed"),
  2201 => (x"c2",x"4b",x"c1",x"87"),
  2202 => (x"c2",x"4b",x"c0",x"87"),
  2203 => (x"c4",x"5b",x"f1",x"d6"),
  2204 => (x"f1",x"d6",x"c2",x"87"),
  2205 => (x"ed",x"d6",x"c2",x"5a"),
  2206 => (x"9a",x"c1",x"4a",x"bf"),
  2207 => (x"49",x"a2",x"c0",x"c1"),
  2208 => (x"fc",x"87",x"e8",x"ec"),
  2209 => (x"ed",x"d6",x"c2",x"48"),
  2210 => (x"ef",x"fe",x"78",x"bf"),
  2211 => (x"4a",x"71",x"1e",x"87"),
  2212 => (x"72",x"1e",x"66",x"c4"),
  2213 => (x"87",x"e2",x"e6",x"49"),
  2214 => (x"1e",x"4f",x"26",x"26"),
  2215 => (x"bf",x"ed",x"d6",x"c2"),
  2216 => (x"87",x"c4",x"e3",x"49"),
  2217 => (x"48",x"c9",x"f1",x"c2"),
  2218 => (x"c2",x"78",x"bf",x"e8"),
  2219 => (x"ec",x"48",x"c5",x"f1"),
  2220 => (x"f1",x"c2",x"78",x"bf"),
  2221 => (x"49",x"4a",x"bf",x"c9"),
  2222 => (x"c8",x"99",x"ff",x"c3"),
  2223 => (x"48",x"72",x"2a",x"b7"),
  2224 => (x"f1",x"c2",x"b0",x"71"),
  2225 => (x"4f",x"26",x"58",x"d1"),
  2226 => (x"5c",x"5b",x"5e",x"0e"),
  2227 => (x"4b",x"71",x"0e",x"5d"),
  2228 => (x"c2",x"87",x"c8",x"ff"),
  2229 => (x"c0",x"48",x"c4",x"f1"),
  2230 => (x"e2",x"49",x"73",x"50"),
  2231 => (x"49",x"70",x"87",x"ea"),
  2232 => (x"cb",x"9c",x"c2",x"4c"),
  2233 => (x"cc",x"cb",x"49",x"ee"),
  2234 => (x"4d",x"49",x"70",x"87"),
  2235 => (x"97",x"c4",x"f1",x"c2"),
  2236 => (x"e2",x"c1",x"05",x"bf"),
  2237 => (x"49",x"66",x"d0",x"87"),
  2238 => (x"bf",x"cd",x"f1",x"c2"),
  2239 => (x"87",x"d6",x"05",x"99"),
  2240 => (x"c2",x"49",x"66",x"d4"),
  2241 => (x"99",x"bf",x"c5",x"f1"),
  2242 => (x"73",x"87",x"cb",x"05"),
  2243 => (x"87",x"f8",x"e1",x"49"),
  2244 => (x"c1",x"02",x"98",x"70"),
  2245 => (x"4c",x"c1",x"87",x"c1"),
  2246 => (x"75",x"87",x"c0",x"fe"),
  2247 => (x"87",x"e1",x"ca",x"49"),
  2248 => (x"c6",x"02",x"98",x"70"),
  2249 => (x"c4",x"f1",x"c2",x"87"),
  2250 => (x"c2",x"50",x"c1",x"48"),
  2251 => (x"bf",x"97",x"c4",x"f1"),
  2252 => (x"87",x"e3",x"c0",x"05"),
  2253 => (x"bf",x"cd",x"f1",x"c2"),
  2254 => (x"99",x"66",x"d0",x"49"),
  2255 => (x"87",x"d6",x"ff",x"05"),
  2256 => (x"bf",x"c5",x"f1",x"c2"),
  2257 => (x"99",x"66",x"d4",x"49"),
  2258 => (x"87",x"ca",x"ff",x"05"),
  2259 => (x"f7",x"e0",x"49",x"73"),
  2260 => (x"05",x"98",x"70",x"87"),
  2261 => (x"74",x"87",x"ff",x"fe"),
  2262 => (x"87",x"dc",x"fb",x"48"),
  2263 => (x"5c",x"5b",x"5e",x"0e"),
  2264 => (x"86",x"f4",x"0e",x"5d"),
  2265 => (x"ec",x"4c",x"4d",x"c0"),
  2266 => (x"a6",x"c4",x"7e",x"bf"),
  2267 => (x"d1",x"f1",x"c2",x"48"),
  2268 => (x"1e",x"c1",x"78",x"bf"),
  2269 => (x"49",x"c7",x"1e",x"c0"),
  2270 => (x"c8",x"87",x"cd",x"fd"),
  2271 => (x"02",x"98",x"70",x"86"),
  2272 => (x"49",x"ff",x"87",x"ce"),
  2273 => (x"c1",x"87",x"cc",x"fb"),
  2274 => (x"df",x"ff",x"49",x"da"),
  2275 => (x"4d",x"c1",x"87",x"fa"),
  2276 => (x"97",x"c4",x"f1",x"c2"),
  2277 => (x"87",x"c3",x"02",x"bf"),
  2278 => (x"c2",x"87",x"c4",x"d0"),
  2279 => (x"4b",x"bf",x"c9",x"f1"),
  2280 => (x"bf",x"ed",x"d6",x"c2"),
  2281 => (x"87",x"eb",x"c0",x"05"),
  2282 => (x"ff",x"49",x"fd",x"c3"),
  2283 => (x"c3",x"87",x"d9",x"df"),
  2284 => (x"df",x"ff",x"49",x"fa"),
  2285 => (x"49",x"73",x"87",x"d2"),
  2286 => (x"71",x"99",x"ff",x"c3"),
  2287 => (x"fb",x"49",x"c0",x"1e"),
  2288 => (x"49",x"73",x"87",x"cb"),
  2289 => (x"71",x"29",x"b7",x"c8"),
  2290 => (x"fa",x"49",x"c1",x"1e"),
  2291 => (x"86",x"c8",x"87",x"ff"),
  2292 => (x"c2",x"87",x"c0",x"c6"),
  2293 => (x"4b",x"bf",x"cd",x"f1"),
  2294 => (x"87",x"dd",x"02",x"9b"),
  2295 => (x"bf",x"e9",x"d6",x"c2"),
  2296 => (x"87",x"dd",x"c7",x"49"),
  2297 => (x"c4",x"05",x"98",x"70"),
  2298 => (x"d2",x"4b",x"c0",x"87"),
  2299 => (x"49",x"e0",x"c2",x"87"),
  2300 => (x"c2",x"87",x"c2",x"c7"),
  2301 => (x"c6",x"58",x"ed",x"d6"),
  2302 => (x"e9",x"d6",x"c2",x"87"),
  2303 => (x"73",x"78",x"c0",x"48"),
  2304 => (x"05",x"99",x"c2",x"49"),
  2305 => (x"eb",x"c3",x"87",x"ce"),
  2306 => (x"fb",x"dd",x"ff",x"49"),
  2307 => (x"c2",x"49",x"70",x"87"),
  2308 => (x"87",x"c2",x"02",x"99"),
  2309 => (x"49",x"73",x"4c",x"fb"),
  2310 => (x"ce",x"05",x"99",x"c1"),
  2311 => (x"49",x"f4",x"c3",x"87"),
  2312 => (x"87",x"e4",x"dd",x"ff"),
  2313 => (x"99",x"c2",x"49",x"70"),
  2314 => (x"fa",x"87",x"c2",x"02"),
  2315 => (x"c8",x"49",x"73",x"4c"),
  2316 => (x"87",x"ce",x"05",x"99"),
  2317 => (x"ff",x"49",x"f5",x"c3"),
  2318 => (x"70",x"87",x"cd",x"dd"),
  2319 => (x"02",x"99",x"c2",x"49"),
  2320 => (x"f1",x"c2",x"87",x"d5"),
  2321 => (x"ca",x"02",x"bf",x"d5"),
  2322 => (x"88",x"c1",x"48",x"87"),
  2323 => (x"58",x"d9",x"f1",x"c2"),
  2324 => (x"ff",x"87",x"c2",x"c0"),
  2325 => (x"73",x"4d",x"c1",x"4c"),
  2326 => (x"05",x"99",x"c4",x"49"),
  2327 => (x"f2",x"c3",x"87",x"ce"),
  2328 => (x"e3",x"dc",x"ff",x"49"),
  2329 => (x"c2",x"49",x"70",x"87"),
  2330 => (x"87",x"dc",x"02",x"99"),
  2331 => (x"bf",x"d5",x"f1",x"c2"),
  2332 => (x"b7",x"c7",x"48",x"7e"),
  2333 => (x"cb",x"c0",x"03",x"a8"),
  2334 => (x"c1",x"48",x"6e",x"87"),
  2335 => (x"d9",x"f1",x"c2",x"80"),
  2336 => (x"87",x"c2",x"c0",x"58"),
  2337 => (x"4d",x"c1",x"4c",x"fe"),
  2338 => (x"ff",x"49",x"fd",x"c3"),
  2339 => (x"70",x"87",x"f9",x"db"),
  2340 => (x"02",x"99",x"c2",x"49"),
  2341 => (x"f1",x"c2",x"87",x"d5"),
  2342 => (x"c0",x"02",x"bf",x"d5"),
  2343 => (x"f1",x"c2",x"87",x"c9"),
  2344 => (x"78",x"c0",x"48",x"d5"),
  2345 => (x"fd",x"87",x"c2",x"c0"),
  2346 => (x"c3",x"4d",x"c1",x"4c"),
  2347 => (x"db",x"ff",x"49",x"fa"),
  2348 => (x"49",x"70",x"87",x"d6"),
  2349 => (x"c0",x"02",x"99",x"c2"),
  2350 => (x"f1",x"c2",x"87",x"d9"),
  2351 => (x"c7",x"48",x"bf",x"d5"),
  2352 => (x"c0",x"03",x"a8",x"b7"),
  2353 => (x"f1",x"c2",x"87",x"c9"),
  2354 => (x"78",x"c7",x"48",x"d5"),
  2355 => (x"fc",x"87",x"c2",x"c0"),
  2356 => (x"c0",x"4d",x"c1",x"4c"),
  2357 => (x"c0",x"03",x"ac",x"b7"),
  2358 => (x"66",x"c4",x"87",x"d1"),
  2359 => (x"82",x"d8",x"c1",x"4a"),
  2360 => (x"c6",x"c0",x"02",x"6a"),
  2361 => (x"74",x"4b",x"6a",x"87"),
  2362 => (x"c0",x"0f",x"73",x"49"),
  2363 => (x"1e",x"f0",x"c3",x"1e"),
  2364 => (x"f7",x"49",x"da",x"c1"),
  2365 => (x"86",x"c8",x"87",x"d2"),
  2366 => (x"c0",x"02",x"98",x"70"),
  2367 => (x"a6",x"c8",x"87",x"e2"),
  2368 => (x"d5",x"f1",x"c2",x"48"),
  2369 => (x"66",x"c8",x"78",x"bf"),
  2370 => (x"c4",x"91",x"cb",x"49"),
  2371 => (x"80",x"71",x"48",x"66"),
  2372 => (x"bf",x"6e",x"7e",x"70"),
  2373 => (x"87",x"c8",x"c0",x"02"),
  2374 => (x"c8",x"4b",x"bf",x"6e"),
  2375 => (x"0f",x"73",x"49",x"66"),
  2376 => (x"c0",x"02",x"9d",x"75"),
  2377 => (x"f1",x"c2",x"87",x"c8"),
  2378 => (x"f3",x"49",x"bf",x"d5"),
  2379 => (x"d6",x"c2",x"87",x"c0"),
  2380 => (x"c0",x"02",x"bf",x"f1"),
  2381 => (x"c2",x"49",x"87",x"dd"),
  2382 => (x"98",x"70",x"87",x"c7"),
  2383 => (x"87",x"d3",x"c0",x"02"),
  2384 => (x"bf",x"d5",x"f1",x"c2"),
  2385 => (x"87",x"e6",x"f2",x"49"),
  2386 => (x"c6",x"f4",x"49",x"c0"),
  2387 => (x"f1",x"d6",x"c2",x"87"),
  2388 => (x"f4",x"78",x"c0",x"48"),
  2389 => (x"87",x"e0",x"f3",x"8e"),
  2390 => (x"5c",x"5b",x"5e",x"0e"),
  2391 => (x"71",x"1e",x"0e",x"5d"),
  2392 => (x"d1",x"f1",x"c2",x"4c"),
  2393 => (x"cd",x"c1",x"49",x"bf"),
  2394 => (x"d1",x"c1",x"4d",x"a1"),
  2395 => (x"74",x"7e",x"69",x"81"),
  2396 => (x"87",x"cf",x"02",x"9c"),
  2397 => (x"74",x"4b",x"a5",x"c4"),
  2398 => (x"d1",x"f1",x"c2",x"7b"),
  2399 => (x"ff",x"f2",x"49",x"bf"),
  2400 => (x"74",x"7b",x"6e",x"87"),
  2401 => (x"87",x"c4",x"05",x"9c"),
  2402 => (x"87",x"c2",x"4b",x"c0"),
  2403 => (x"49",x"73",x"4b",x"c1"),
  2404 => (x"d4",x"87",x"c0",x"f3"),
  2405 => (x"87",x"c7",x"02",x"66"),
  2406 => (x"70",x"87",x"da",x"49"),
  2407 => (x"c0",x"87",x"c2",x"4a"),
  2408 => (x"f5",x"d6",x"c2",x"4a"),
  2409 => (x"cf",x"f2",x"26",x"5a"),
  2410 => (x"00",x"00",x"00",x"87"),
  2411 => (x"00",x"00",x"00",x"00"),
  2412 => (x"00",x"00",x"00",x"00"),
  2413 => (x"4a",x"71",x"1e",x"00"),
  2414 => (x"49",x"bf",x"c8",x"ff"),
  2415 => (x"26",x"48",x"a1",x"72"),
  2416 => (x"c8",x"ff",x"1e",x"4f"),
  2417 => (x"c0",x"fe",x"89",x"bf"),
  2418 => (x"c0",x"c0",x"c0",x"c0"),
  2419 => (x"87",x"c4",x"01",x"a9"),
  2420 => (x"87",x"c2",x"4a",x"c0"),
  2421 => (x"48",x"72",x"4a",x"c1"),
  2422 => (x"5e",x"0e",x"4f",x"26"),
  2423 => (x"0e",x"5d",x"5c",x"5b"),
  2424 => (x"d4",x"ff",x"4b",x"71"),
  2425 => (x"48",x"66",x"d0",x"4c"),
  2426 => (x"49",x"d6",x"78",x"c0"),
  2427 => (x"87",x"d0",x"d8",x"ff"),
  2428 => (x"6c",x"7c",x"ff",x"c3"),
  2429 => (x"99",x"ff",x"c3",x"49"),
  2430 => (x"c3",x"49",x"4d",x"71"),
  2431 => (x"e0",x"c1",x"99",x"f0"),
  2432 => (x"87",x"cb",x"05",x"a9"),
  2433 => (x"6c",x"7c",x"ff",x"c3"),
  2434 => (x"d0",x"98",x"c3",x"48"),
  2435 => (x"c3",x"78",x"08",x"66"),
  2436 => (x"4a",x"6c",x"7c",x"ff"),
  2437 => (x"c3",x"31",x"c8",x"49"),
  2438 => (x"4a",x"6c",x"7c",x"ff"),
  2439 => (x"49",x"72",x"b2",x"71"),
  2440 => (x"ff",x"c3",x"31",x"c8"),
  2441 => (x"71",x"4a",x"6c",x"7c"),
  2442 => (x"c8",x"49",x"72",x"b2"),
  2443 => (x"7c",x"ff",x"c3",x"31"),
  2444 => (x"b2",x"71",x"4a",x"6c"),
  2445 => (x"c0",x"48",x"d0",x"ff"),
  2446 => (x"9b",x"73",x"78",x"e0"),
  2447 => (x"72",x"87",x"c2",x"02"),
  2448 => (x"26",x"48",x"75",x"7b"),
  2449 => (x"26",x"4c",x"26",x"4d"),
  2450 => (x"1e",x"4f",x"26",x"4b"),
  2451 => (x"5e",x"0e",x"4f",x"26"),
  2452 => (x"f8",x"0e",x"5c",x"5b"),
  2453 => (x"c8",x"1e",x"76",x"86"),
  2454 => (x"fd",x"fd",x"49",x"a6"),
  2455 => (x"70",x"86",x"c4",x"87"),
  2456 => (x"c2",x"48",x"6e",x"4b"),
  2457 => (x"f0",x"c2",x"03",x"a8"),
  2458 => (x"c3",x"4a",x"73",x"87"),
  2459 => (x"d0",x"c1",x"9a",x"f0"),
  2460 => (x"87",x"c7",x"02",x"aa"),
  2461 => (x"05",x"aa",x"e0",x"c1"),
  2462 => (x"73",x"87",x"de",x"c2"),
  2463 => (x"02",x"99",x"c8",x"49"),
  2464 => (x"c6",x"ff",x"87",x"c3"),
  2465 => (x"c3",x"4c",x"73",x"87"),
  2466 => (x"05",x"ac",x"c2",x"9c"),
  2467 => (x"c4",x"87",x"c2",x"c1"),
  2468 => (x"31",x"c9",x"49",x"66"),
  2469 => (x"66",x"c4",x"1e",x"71"),
  2470 => (x"c2",x"92",x"d4",x"4a"),
  2471 => (x"72",x"49",x"d9",x"f1"),
  2472 => (x"ed",x"cc",x"fe",x"81"),
  2473 => (x"ff",x"49",x"d8",x"87"),
  2474 => (x"c8",x"87",x"d5",x"d5"),
  2475 => (x"df",x"c2",x"1e",x"c0"),
  2476 => (x"e8",x"fd",x"49",x"f2"),
  2477 => (x"d0",x"ff",x"87",x"e9"),
  2478 => (x"78",x"e0",x"c0",x"48"),
  2479 => (x"1e",x"f2",x"df",x"c2"),
  2480 => (x"d4",x"4a",x"66",x"cc"),
  2481 => (x"d9",x"f1",x"c2",x"92"),
  2482 => (x"fe",x"81",x"72",x"49"),
  2483 => (x"cc",x"87",x"f4",x"ca"),
  2484 => (x"05",x"ac",x"c1",x"86"),
  2485 => (x"c4",x"87",x"c2",x"c1"),
  2486 => (x"31",x"c9",x"49",x"66"),
  2487 => (x"66",x"c4",x"1e",x"71"),
  2488 => (x"c2",x"92",x"d4",x"4a"),
  2489 => (x"72",x"49",x"d9",x"f1"),
  2490 => (x"e5",x"cb",x"fe",x"81"),
  2491 => (x"f2",x"df",x"c2",x"87"),
  2492 => (x"4a",x"66",x"c8",x"1e"),
  2493 => (x"f1",x"c2",x"92",x"d4"),
  2494 => (x"81",x"72",x"49",x"d9"),
  2495 => (x"87",x"f4",x"c8",x"fe"),
  2496 => (x"d3",x"ff",x"49",x"d7"),
  2497 => (x"c0",x"c8",x"87",x"fa"),
  2498 => (x"f2",x"df",x"c2",x"1e"),
  2499 => (x"e7",x"e6",x"fd",x"49"),
  2500 => (x"ff",x"86",x"cc",x"87"),
  2501 => (x"e0",x"c0",x"48",x"d0"),
  2502 => (x"fc",x"8e",x"f8",x"78"),
  2503 => (x"5e",x"0e",x"87",x"e7"),
  2504 => (x"0e",x"5d",x"5c",x"5b"),
  2505 => (x"ff",x"4d",x"71",x"1e"),
  2506 => (x"66",x"d4",x"4c",x"d4"),
  2507 => (x"b7",x"c3",x"48",x"7e"),
  2508 => (x"87",x"c5",x"06",x"a8"),
  2509 => (x"e2",x"c1",x"48",x"c0"),
  2510 => (x"fe",x"49",x"75",x"87"),
  2511 => (x"75",x"87",x"f8",x"d9"),
  2512 => (x"4b",x"66",x"c4",x"1e"),
  2513 => (x"f1",x"c2",x"93",x"d4"),
  2514 => (x"49",x"73",x"83",x"d9"),
  2515 => (x"87",x"f1",x"c2",x"fe"),
  2516 => (x"4b",x"6b",x"83",x"c8"),
  2517 => (x"c8",x"48",x"d0",x"ff"),
  2518 => (x"7c",x"dd",x"78",x"e1"),
  2519 => (x"ff",x"c3",x"49",x"73"),
  2520 => (x"73",x"7c",x"71",x"99"),
  2521 => (x"29",x"b7",x"c8",x"49"),
  2522 => (x"71",x"99",x"ff",x"c3"),
  2523 => (x"d0",x"49",x"73",x"7c"),
  2524 => (x"ff",x"c3",x"29",x"b7"),
  2525 => (x"73",x"7c",x"71",x"99"),
  2526 => (x"29",x"b7",x"d8",x"49"),
  2527 => (x"7c",x"c0",x"7c",x"71"),
  2528 => (x"7c",x"7c",x"7c",x"7c"),
  2529 => (x"7c",x"7c",x"7c",x"7c"),
  2530 => (x"c0",x"7c",x"7c",x"7c"),
  2531 => (x"66",x"c4",x"78",x"e0"),
  2532 => (x"ff",x"49",x"dc",x"1e"),
  2533 => (x"c8",x"87",x"ce",x"d2"),
  2534 => (x"26",x"48",x"73",x"86"),
  2535 => (x"1e",x"87",x"e4",x"fa"),
  2536 => (x"bf",x"c8",x"df",x"c2"),
  2537 => (x"c2",x"b9",x"c1",x"49"),
  2538 => (x"ff",x"59",x"cc",x"df"),
  2539 => (x"ff",x"c3",x"48",x"d4"),
  2540 => (x"48",x"d0",x"ff",x"78"),
  2541 => (x"ff",x"78",x"e1",x"c0"),
  2542 => (x"78",x"c1",x"48",x"d4"),
  2543 => (x"78",x"71",x"31",x"c4"),
  2544 => (x"c0",x"48",x"d0",x"ff"),
  2545 => (x"4f",x"26",x"78",x"e0"),
  2546 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

