package build_id is
constant BUILD_DATE : string := "230418";
constant BUILD_TIME : string := "211450";
end build_id;
