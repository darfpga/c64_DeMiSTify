package build_id is
constant BUILD_DATE : string := "230331";
constant BUILD_TIME : string := "133318";
end build_id;
