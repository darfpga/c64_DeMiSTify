
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f0",x"f1",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"f0",x"f1",x"c2"),
    14 => (x"48",x"f8",x"de",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"d9",x"e1"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"4a",x"71",x"1e",x"4f"),
    50 => (x"48",x"49",x"66",x"c4"),
    51 => (x"a6",x"c8",x"88",x"c1"),
    52 => (x"02",x"99",x"71",x"58"),
    53 => (x"48",x"12",x"87",x"d4"),
    54 => (x"78",x"08",x"d4",x"ff"),
    55 => (x"48",x"49",x"66",x"c4"),
    56 => (x"a6",x"c8",x"88",x"c1"),
    57 => (x"05",x"99",x"71",x"58"),
    58 => (x"4f",x"26",x"87",x"ec"),
    59 => (x"c4",x"4a",x"71",x"1e"),
    60 => (x"c1",x"48",x"49",x"66"),
    61 => (x"58",x"a6",x"c8",x"88"),
    62 => (x"d6",x"02",x"99",x"71"),
    63 => (x"48",x"d4",x"ff",x"87"),
    64 => (x"68",x"78",x"ff",x"c3"),
    65 => (x"49",x"66",x"c4",x"52"),
    66 => (x"c8",x"88",x"c1",x"48"),
    67 => (x"99",x"71",x"58",x"a6"),
    68 => (x"26",x"87",x"ea",x"05"),
    69 => (x"1e",x"73",x"1e",x"4f"),
    70 => (x"c3",x"4b",x"d4",x"ff"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"6b",x"7b",x"ff",x"c3"),
    73 => (x"72",x"32",x"c8",x"49"),
    74 => (x"7b",x"ff",x"c3",x"b1"),
    75 => (x"31",x"c8",x"4a",x"6b"),
    76 => (x"ff",x"c3",x"b2",x"71"),
    77 => (x"c8",x"49",x"6b",x"7b"),
    78 => (x"71",x"b1",x"72",x"32"),
    79 => (x"26",x"87",x"c4",x"48"),
    80 => (x"26",x"4c",x"26",x"4d"),
    81 => (x"0e",x"4f",x"26",x"4b"),
    82 => (x"5d",x"5c",x"5b",x"5e"),
    83 => (x"ff",x"4a",x"71",x"0e"),
    84 => (x"49",x"72",x"4c",x"d4"),
    85 => (x"71",x"99",x"ff",x"c3"),
    86 => (x"f8",x"de",x"c2",x"7c"),
    87 => (x"87",x"c8",x"05",x"bf"),
    88 => (x"c9",x"48",x"66",x"d0"),
    89 => (x"58",x"a6",x"d4",x"30"),
    90 => (x"d8",x"49",x"66",x"d0"),
    91 => (x"99",x"ff",x"c3",x"29"),
    92 => (x"66",x"d0",x"7c",x"71"),
    93 => (x"c3",x"29",x"d0",x"49"),
    94 => (x"7c",x"71",x"99",x"ff"),
    95 => (x"c8",x"49",x"66",x"d0"),
    96 => (x"99",x"ff",x"c3",x"29"),
    97 => (x"66",x"d0",x"7c",x"71"),
    98 => (x"99",x"ff",x"c3",x"49"),
    99 => (x"49",x"72",x"7c",x"71"),
   100 => (x"ff",x"c3",x"29",x"d0"),
   101 => (x"6c",x"7c",x"71",x"99"),
   102 => (x"ff",x"f0",x"c9",x"4b"),
   103 => (x"ab",x"ff",x"c3",x"4d"),
   104 => (x"c3",x"87",x"d0",x"05"),
   105 => (x"4b",x"6c",x"7c",x"ff"),
   106 => (x"c6",x"02",x"8d",x"c1"),
   107 => (x"ab",x"ff",x"c3",x"87"),
   108 => (x"73",x"87",x"f0",x"02"),
   109 => (x"87",x"c7",x"fe",x"48"),
   110 => (x"ff",x"49",x"c0",x"1e"),
   111 => (x"ff",x"c3",x"48",x"d4"),
   112 => (x"c3",x"81",x"c1",x"78"),
   113 => (x"04",x"a9",x"b7",x"c8"),
   114 => (x"4f",x"26",x"87",x"f1"),
   115 => (x"e7",x"1e",x"73",x"1e"),
   116 => (x"df",x"f8",x"c4",x"87"),
   117 => (x"c0",x"1e",x"c0",x"4b"),
   118 => (x"f7",x"c1",x"f0",x"ff"),
   119 => (x"87",x"e7",x"fd",x"49"),
   120 => (x"a8",x"c1",x"86",x"c4"),
   121 => (x"87",x"ea",x"c0",x"05"),
   122 => (x"c3",x"48",x"d4",x"ff"),
   123 => (x"c0",x"c1",x"78",x"ff"),
   124 => (x"c0",x"c0",x"c0",x"c0"),
   125 => (x"f0",x"e1",x"c0",x"1e"),
   126 => (x"fd",x"49",x"e9",x"c1"),
   127 => (x"86",x"c4",x"87",x"c9"),
   128 => (x"ca",x"05",x"98",x"70"),
   129 => (x"48",x"d4",x"ff",x"87"),
   130 => (x"c1",x"78",x"ff",x"c3"),
   131 => (x"fe",x"87",x"cb",x"48"),
   132 => (x"8b",x"c1",x"87",x"e6"),
   133 => (x"87",x"fd",x"fe",x"05"),
   134 => (x"e6",x"fc",x"48",x"c0"),
   135 => (x"1e",x"73",x"1e",x"87"),
   136 => (x"c3",x"48",x"d4",x"ff"),
   137 => (x"4b",x"d3",x"78",x"ff"),
   138 => (x"ff",x"c0",x"1e",x"c0"),
   139 => (x"49",x"c1",x"c1",x"f0"),
   140 => (x"c4",x"87",x"d4",x"fc"),
   141 => (x"05",x"98",x"70",x"86"),
   142 => (x"d4",x"ff",x"87",x"ca"),
   143 => (x"78",x"ff",x"c3",x"48"),
   144 => (x"87",x"cb",x"48",x"c1"),
   145 => (x"c1",x"87",x"f1",x"fd"),
   146 => (x"db",x"ff",x"05",x"8b"),
   147 => (x"fb",x"48",x"c0",x"87"),
   148 => (x"5e",x"0e",x"87",x"f1"),
   149 => (x"ff",x"0e",x"5c",x"5b"),
   150 => (x"db",x"fd",x"4c",x"d4"),
   151 => (x"1e",x"ea",x"c6",x"87"),
   152 => (x"c1",x"f0",x"e1",x"c0"),
   153 => (x"de",x"fb",x"49",x"c8"),
   154 => (x"c1",x"86",x"c4",x"87"),
   155 => (x"87",x"c8",x"02",x"a8"),
   156 => (x"c0",x"87",x"ea",x"fe"),
   157 => (x"87",x"e2",x"c1",x"48"),
   158 => (x"70",x"87",x"da",x"fa"),
   159 => (x"ff",x"ff",x"cf",x"49"),
   160 => (x"a9",x"ea",x"c6",x"99"),
   161 => (x"fe",x"87",x"c8",x"02"),
   162 => (x"48",x"c0",x"87",x"d3"),
   163 => (x"c3",x"87",x"cb",x"c1"),
   164 => (x"f1",x"c0",x"7c",x"ff"),
   165 => (x"87",x"f4",x"fc",x"4b"),
   166 => (x"c0",x"02",x"98",x"70"),
   167 => (x"1e",x"c0",x"87",x"eb"),
   168 => (x"c1",x"f0",x"ff",x"c0"),
   169 => (x"de",x"fa",x"49",x"fa"),
   170 => (x"70",x"86",x"c4",x"87"),
   171 => (x"87",x"d9",x"05",x"98"),
   172 => (x"6c",x"7c",x"ff",x"c3"),
   173 => (x"7c",x"ff",x"c3",x"49"),
   174 => (x"c1",x"7c",x"7c",x"7c"),
   175 => (x"c4",x"02",x"99",x"c0"),
   176 => (x"d5",x"48",x"c1",x"87"),
   177 => (x"d1",x"48",x"c0",x"87"),
   178 => (x"05",x"ab",x"c2",x"87"),
   179 => (x"48",x"c0",x"87",x"c4"),
   180 => (x"8b",x"c1",x"87",x"c8"),
   181 => (x"87",x"fd",x"fe",x"05"),
   182 => (x"e4",x"f9",x"48",x"c0"),
   183 => (x"1e",x"73",x"1e",x"87"),
   184 => (x"48",x"f8",x"de",x"c2"),
   185 => (x"4b",x"c7",x"78",x"c1"),
   186 => (x"c2",x"48",x"d0",x"ff"),
   187 => (x"87",x"c8",x"fb",x"78"),
   188 => (x"c3",x"48",x"d0",x"ff"),
   189 => (x"c0",x"1e",x"c0",x"78"),
   190 => (x"c0",x"c1",x"d0",x"e5"),
   191 => (x"87",x"c7",x"f9",x"49"),
   192 => (x"a8",x"c1",x"86",x"c4"),
   193 => (x"4b",x"87",x"c1",x"05"),
   194 => (x"c5",x"05",x"ab",x"c2"),
   195 => (x"c0",x"48",x"c0",x"87"),
   196 => (x"8b",x"c1",x"87",x"f9"),
   197 => (x"87",x"d0",x"ff",x"05"),
   198 => (x"c2",x"87",x"f7",x"fc"),
   199 => (x"70",x"58",x"fc",x"de"),
   200 => (x"87",x"cd",x"05",x"98"),
   201 => (x"ff",x"c0",x"1e",x"c1"),
   202 => (x"49",x"d0",x"c1",x"f0"),
   203 => (x"c4",x"87",x"d8",x"f8"),
   204 => (x"48",x"d4",x"ff",x"86"),
   205 => (x"c4",x"78",x"ff",x"c3"),
   206 => (x"df",x"c2",x"87",x"de"),
   207 => (x"d0",x"ff",x"58",x"c0"),
   208 => (x"ff",x"78",x"c2",x"48"),
   209 => (x"ff",x"c3",x"48",x"d4"),
   210 => (x"f7",x"48",x"c1",x"78"),
   211 => (x"5e",x"0e",x"87",x"f5"),
   212 => (x"0e",x"5d",x"5c",x"5b"),
   213 => (x"ff",x"c3",x"4a",x"71"),
   214 => (x"4c",x"d4",x"ff",x"4d"),
   215 => (x"d0",x"ff",x"7c",x"75"),
   216 => (x"78",x"c3",x"c4",x"48"),
   217 => (x"1e",x"72",x"7c",x"75"),
   218 => (x"c1",x"f0",x"ff",x"c0"),
   219 => (x"d6",x"f7",x"49",x"d8"),
   220 => (x"70",x"86",x"c4",x"87"),
   221 => (x"87",x"c5",x"02",x"98"),
   222 => (x"f0",x"c0",x"48",x"c1"),
   223 => (x"c3",x"7c",x"75",x"87"),
   224 => (x"c0",x"c8",x"7c",x"fe"),
   225 => (x"49",x"66",x"d4",x"1e"),
   226 => (x"c4",x"87",x"fa",x"f4"),
   227 => (x"75",x"7c",x"75",x"86"),
   228 => (x"d8",x"7c",x"75",x"7c"),
   229 => (x"75",x"4b",x"e0",x"da"),
   230 => (x"99",x"49",x"6c",x"7c"),
   231 => (x"c1",x"87",x"c5",x"05"),
   232 => (x"87",x"f3",x"05",x"8b"),
   233 => (x"d0",x"ff",x"7c",x"75"),
   234 => (x"c0",x"78",x"c2",x"48"),
   235 => (x"87",x"cf",x"f6",x"48"),
   236 => (x"5c",x"5b",x"5e",x"0e"),
   237 => (x"4b",x"71",x"0e",x"5d"),
   238 => (x"ee",x"c5",x"4c",x"c0"),
   239 => (x"ff",x"4a",x"df",x"cd"),
   240 => (x"ff",x"c3",x"48",x"d4"),
   241 => (x"c3",x"49",x"68",x"78"),
   242 => (x"c0",x"05",x"a9",x"fe"),
   243 => (x"4d",x"70",x"87",x"fd"),
   244 => (x"cc",x"02",x"9b",x"73"),
   245 => (x"1e",x"66",x"d0",x"87"),
   246 => (x"cf",x"f4",x"49",x"73"),
   247 => (x"d6",x"86",x"c4",x"87"),
   248 => (x"48",x"d0",x"ff",x"87"),
   249 => (x"c3",x"78",x"d1",x"c4"),
   250 => (x"66",x"d0",x"7d",x"ff"),
   251 => (x"d4",x"88",x"c1",x"48"),
   252 => (x"98",x"70",x"58",x"a6"),
   253 => (x"ff",x"87",x"f0",x"05"),
   254 => (x"ff",x"c3",x"48",x"d4"),
   255 => (x"9b",x"73",x"78",x"78"),
   256 => (x"ff",x"87",x"c5",x"05"),
   257 => (x"78",x"d0",x"48",x"d0"),
   258 => (x"c1",x"4c",x"4a",x"c1"),
   259 => (x"ee",x"fe",x"05",x"8a"),
   260 => (x"f4",x"48",x"74",x"87"),
   261 => (x"73",x"1e",x"87",x"e9"),
   262 => (x"c0",x"4a",x"71",x"1e"),
   263 => (x"48",x"d4",x"ff",x"4b"),
   264 => (x"ff",x"78",x"ff",x"c3"),
   265 => (x"c3",x"c4",x"48",x"d0"),
   266 => (x"48",x"d4",x"ff",x"78"),
   267 => (x"72",x"78",x"ff",x"c3"),
   268 => (x"f0",x"ff",x"c0",x"1e"),
   269 => (x"f4",x"49",x"d1",x"c1"),
   270 => (x"86",x"c4",x"87",x"cd"),
   271 => (x"d2",x"05",x"98",x"70"),
   272 => (x"1e",x"c0",x"c8",x"87"),
   273 => (x"fd",x"49",x"66",x"cc"),
   274 => (x"86",x"c4",x"87",x"e6"),
   275 => (x"d0",x"ff",x"4b",x"70"),
   276 => (x"73",x"78",x"c2",x"48"),
   277 => (x"87",x"eb",x"f3",x"48"),
   278 => (x"5c",x"5b",x"5e",x"0e"),
   279 => (x"1e",x"c0",x"0e",x"5d"),
   280 => (x"c1",x"f0",x"ff",x"c0"),
   281 => (x"de",x"f3",x"49",x"c9"),
   282 => (x"c2",x"1e",x"d2",x"87"),
   283 => (x"fc",x"49",x"c0",x"df"),
   284 => (x"86",x"c8",x"87",x"fe"),
   285 => (x"84",x"c1",x"4c",x"c0"),
   286 => (x"04",x"ac",x"b7",x"d2"),
   287 => (x"df",x"c2",x"87",x"f8"),
   288 => (x"49",x"bf",x"97",x"c0"),
   289 => (x"c1",x"99",x"c0",x"c3"),
   290 => (x"c0",x"05",x"a9",x"c0"),
   291 => (x"df",x"c2",x"87",x"e7"),
   292 => (x"49",x"bf",x"97",x"c7"),
   293 => (x"df",x"c2",x"31",x"d0"),
   294 => (x"4a",x"bf",x"97",x"c8"),
   295 => (x"b1",x"72",x"32",x"c8"),
   296 => (x"97",x"c9",x"df",x"c2"),
   297 => (x"71",x"b1",x"4a",x"bf"),
   298 => (x"ff",x"ff",x"cf",x"4c"),
   299 => (x"84",x"c1",x"9c",x"ff"),
   300 => (x"e7",x"c1",x"34",x"ca"),
   301 => (x"c9",x"df",x"c2",x"87"),
   302 => (x"c1",x"49",x"bf",x"97"),
   303 => (x"c2",x"99",x"c6",x"31"),
   304 => (x"bf",x"97",x"ca",x"df"),
   305 => (x"2a",x"b7",x"c7",x"4a"),
   306 => (x"df",x"c2",x"b1",x"72"),
   307 => (x"4a",x"bf",x"97",x"c5"),
   308 => (x"c2",x"9d",x"cf",x"4d"),
   309 => (x"bf",x"97",x"c6",x"df"),
   310 => (x"ca",x"9a",x"c3",x"4a"),
   311 => (x"c7",x"df",x"c2",x"32"),
   312 => (x"c2",x"4b",x"bf",x"97"),
   313 => (x"c2",x"b2",x"73",x"33"),
   314 => (x"bf",x"97",x"c8",x"df"),
   315 => (x"9b",x"c0",x"c3",x"4b"),
   316 => (x"73",x"2b",x"b7",x"c6"),
   317 => (x"c1",x"81",x"c2",x"b2"),
   318 => (x"70",x"30",x"71",x"48"),
   319 => (x"75",x"48",x"c1",x"49"),
   320 => (x"72",x"4d",x"70",x"30"),
   321 => (x"71",x"84",x"c1",x"4c"),
   322 => (x"b7",x"c0",x"c8",x"94"),
   323 => (x"87",x"cc",x"06",x"ad"),
   324 => (x"2d",x"b7",x"34",x"c1"),
   325 => (x"ad",x"b7",x"c0",x"c8"),
   326 => (x"87",x"f4",x"ff",x"01"),
   327 => (x"de",x"f0",x"48",x"74"),
   328 => (x"5b",x"5e",x"0e",x"87"),
   329 => (x"f8",x"0e",x"5d",x"5c"),
   330 => (x"e6",x"e7",x"c2",x"86"),
   331 => (x"c2",x"78",x"c0",x"48"),
   332 => (x"c0",x"1e",x"de",x"df"),
   333 => (x"87",x"de",x"fb",x"49"),
   334 => (x"98",x"70",x"86",x"c4"),
   335 => (x"c0",x"87",x"c5",x"05"),
   336 => (x"87",x"ce",x"c9",x"48"),
   337 => (x"7e",x"c1",x"4d",x"c0"),
   338 => (x"bf",x"c0",x"f3",x"c0"),
   339 => (x"d4",x"e0",x"c2",x"49"),
   340 => (x"4b",x"c8",x"71",x"4a"),
   341 => (x"70",x"87",x"d3",x"ec"),
   342 => (x"87",x"c2",x"05",x"98"),
   343 => (x"f2",x"c0",x"7e",x"c0"),
   344 => (x"c2",x"49",x"bf",x"fc"),
   345 => (x"71",x"4a",x"f0",x"e0"),
   346 => (x"fd",x"eb",x"4b",x"c8"),
   347 => (x"05",x"98",x"70",x"87"),
   348 => (x"7e",x"c0",x"87",x"c2"),
   349 => (x"fd",x"c0",x"02",x"6e"),
   350 => (x"e4",x"e6",x"c2",x"87"),
   351 => (x"e7",x"c2",x"4d",x"bf"),
   352 => (x"7e",x"bf",x"9f",x"dc"),
   353 => (x"ea",x"d6",x"c5",x"48"),
   354 => (x"87",x"c7",x"05",x"a8"),
   355 => (x"bf",x"e4",x"e6",x"c2"),
   356 => (x"6e",x"87",x"ce",x"4d"),
   357 => (x"d5",x"e9",x"ca",x"48"),
   358 => (x"87",x"c5",x"02",x"a8"),
   359 => (x"f1",x"c7",x"48",x"c0"),
   360 => (x"de",x"df",x"c2",x"87"),
   361 => (x"f9",x"49",x"75",x"1e"),
   362 => (x"86",x"c4",x"87",x"ec"),
   363 => (x"c5",x"05",x"98",x"70"),
   364 => (x"c7",x"48",x"c0",x"87"),
   365 => (x"f2",x"c0",x"87",x"dc"),
   366 => (x"c2",x"49",x"bf",x"fc"),
   367 => (x"71",x"4a",x"f0",x"e0"),
   368 => (x"e5",x"ea",x"4b",x"c8"),
   369 => (x"05",x"98",x"70",x"87"),
   370 => (x"e7",x"c2",x"87",x"c8"),
   371 => (x"78",x"c1",x"48",x"e6"),
   372 => (x"f3",x"c0",x"87",x"da"),
   373 => (x"c2",x"49",x"bf",x"c0"),
   374 => (x"71",x"4a",x"d4",x"e0"),
   375 => (x"c9",x"ea",x"4b",x"c8"),
   376 => (x"02",x"98",x"70",x"87"),
   377 => (x"c0",x"87",x"c5",x"c0"),
   378 => (x"87",x"e6",x"c6",x"48"),
   379 => (x"97",x"dc",x"e7",x"c2"),
   380 => (x"d5",x"c1",x"49",x"bf"),
   381 => (x"cd",x"c0",x"05",x"a9"),
   382 => (x"dd",x"e7",x"c2",x"87"),
   383 => (x"c2",x"49",x"bf",x"97"),
   384 => (x"c0",x"02",x"a9",x"ea"),
   385 => (x"48",x"c0",x"87",x"c5"),
   386 => (x"c2",x"87",x"c7",x"c6"),
   387 => (x"bf",x"97",x"de",x"df"),
   388 => (x"e9",x"c3",x"48",x"7e"),
   389 => (x"ce",x"c0",x"02",x"a8"),
   390 => (x"c3",x"48",x"6e",x"87"),
   391 => (x"c0",x"02",x"a8",x"eb"),
   392 => (x"48",x"c0",x"87",x"c5"),
   393 => (x"c2",x"87",x"eb",x"c5"),
   394 => (x"bf",x"97",x"e9",x"df"),
   395 => (x"c0",x"05",x"99",x"49"),
   396 => (x"df",x"c2",x"87",x"cc"),
   397 => (x"49",x"bf",x"97",x"ea"),
   398 => (x"c0",x"02",x"a9",x"c2"),
   399 => (x"48",x"c0",x"87",x"c5"),
   400 => (x"c2",x"87",x"cf",x"c5"),
   401 => (x"bf",x"97",x"eb",x"df"),
   402 => (x"e2",x"e7",x"c2",x"48"),
   403 => (x"48",x"4c",x"70",x"58"),
   404 => (x"e7",x"c2",x"88",x"c1"),
   405 => (x"df",x"c2",x"58",x"e6"),
   406 => (x"49",x"bf",x"97",x"ec"),
   407 => (x"df",x"c2",x"81",x"75"),
   408 => (x"4a",x"bf",x"97",x"ed"),
   409 => (x"a1",x"72",x"32",x"c8"),
   410 => (x"f3",x"eb",x"c2",x"7e"),
   411 => (x"c2",x"78",x"6e",x"48"),
   412 => (x"bf",x"97",x"ee",x"df"),
   413 => (x"58",x"a6",x"c8",x"48"),
   414 => (x"bf",x"e6",x"e7",x"c2"),
   415 => (x"87",x"d4",x"c2",x"02"),
   416 => (x"bf",x"fc",x"f2",x"c0"),
   417 => (x"f0",x"e0",x"c2",x"49"),
   418 => (x"4b",x"c8",x"71",x"4a"),
   419 => (x"70",x"87",x"db",x"e7"),
   420 => (x"c5",x"c0",x"02",x"98"),
   421 => (x"c3",x"48",x"c0",x"87"),
   422 => (x"e7",x"c2",x"87",x"f8"),
   423 => (x"c2",x"4c",x"bf",x"de"),
   424 => (x"c2",x"5c",x"c7",x"ec"),
   425 => (x"bf",x"97",x"c3",x"e0"),
   426 => (x"c2",x"31",x"c8",x"49"),
   427 => (x"bf",x"97",x"c2",x"e0"),
   428 => (x"c2",x"49",x"a1",x"4a"),
   429 => (x"bf",x"97",x"c4",x"e0"),
   430 => (x"72",x"32",x"d0",x"4a"),
   431 => (x"e0",x"c2",x"49",x"a1"),
   432 => (x"4a",x"bf",x"97",x"c5"),
   433 => (x"a1",x"72",x"32",x"d8"),
   434 => (x"91",x"66",x"c4",x"49"),
   435 => (x"bf",x"f3",x"eb",x"c2"),
   436 => (x"fb",x"eb",x"c2",x"81"),
   437 => (x"cb",x"e0",x"c2",x"59"),
   438 => (x"c8",x"4a",x"bf",x"97"),
   439 => (x"ca",x"e0",x"c2",x"32"),
   440 => (x"a2",x"4b",x"bf",x"97"),
   441 => (x"cc",x"e0",x"c2",x"4a"),
   442 => (x"d0",x"4b",x"bf",x"97"),
   443 => (x"4a",x"a2",x"73",x"33"),
   444 => (x"97",x"cd",x"e0",x"c2"),
   445 => (x"9b",x"cf",x"4b",x"bf"),
   446 => (x"a2",x"73",x"33",x"d8"),
   447 => (x"ff",x"eb",x"c2",x"4a"),
   448 => (x"fb",x"eb",x"c2",x"5a"),
   449 => (x"8a",x"c2",x"4a",x"bf"),
   450 => (x"eb",x"c2",x"92",x"74"),
   451 => (x"a1",x"72",x"48",x"ff"),
   452 => (x"87",x"ca",x"c1",x"78"),
   453 => (x"97",x"f0",x"df",x"c2"),
   454 => (x"31",x"c8",x"49",x"bf"),
   455 => (x"97",x"ef",x"df",x"c2"),
   456 => (x"49",x"a1",x"4a",x"bf"),
   457 => (x"59",x"ee",x"e7",x"c2"),
   458 => (x"bf",x"ea",x"e7",x"c2"),
   459 => (x"c7",x"31",x"c5",x"49"),
   460 => (x"29",x"c9",x"81",x"ff"),
   461 => (x"59",x"c7",x"ec",x"c2"),
   462 => (x"97",x"f5",x"df",x"c2"),
   463 => (x"32",x"c8",x"4a",x"bf"),
   464 => (x"97",x"f4",x"df",x"c2"),
   465 => (x"4a",x"a2",x"4b",x"bf"),
   466 => (x"6e",x"92",x"66",x"c4"),
   467 => (x"c3",x"ec",x"c2",x"82"),
   468 => (x"fb",x"eb",x"c2",x"5a"),
   469 => (x"c2",x"78",x"c0",x"48"),
   470 => (x"72",x"48",x"f7",x"eb"),
   471 => (x"ec",x"c2",x"78",x"a1"),
   472 => (x"eb",x"c2",x"48",x"c7"),
   473 => (x"c2",x"78",x"bf",x"fb"),
   474 => (x"c2",x"48",x"cb",x"ec"),
   475 => (x"78",x"bf",x"ff",x"eb"),
   476 => (x"bf",x"e6",x"e7",x"c2"),
   477 => (x"87",x"c9",x"c0",x"02"),
   478 => (x"30",x"c4",x"48",x"74"),
   479 => (x"c9",x"c0",x"7e",x"70"),
   480 => (x"c3",x"ec",x"c2",x"87"),
   481 => (x"30",x"c4",x"48",x"bf"),
   482 => (x"e7",x"c2",x"7e",x"70"),
   483 => (x"78",x"6e",x"48",x"ea"),
   484 => (x"8e",x"f8",x"48",x"c1"),
   485 => (x"4c",x"26",x"4d",x"26"),
   486 => (x"4f",x"26",x"4b",x"26"),
   487 => (x"5c",x"5b",x"5e",x"0e"),
   488 => (x"4a",x"71",x"0e",x"5d"),
   489 => (x"bf",x"e6",x"e7",x"c2"),
   490 => (x"72",x"87",x"cb",x"02"),
   491 => (x"72",x"2b",x"c7",x"4b"),
   492 => (x"9c",x"ff",x"c1",x"4c"),
   493 => (x"4b",x"72",x"87",x"c9"),
   494 => (x"4c",x"72",x"2b",x"c8"),
   495 => (x"c2",x"9c",x"ff",x"c3"),
   496 => (x"83",x"bf",x"f3",x"eb"),
   497 => (x"bf",x"f8",x"f2",x"c0"),
   498 => (x"87",x"d9",x"02",x"ab"),
   499 => (x"5b",x"fc",x"f2",x"c0"),
   500 => (x"1e",x"de",x"df",x"c2"),
   501 => (x"fd",x"f0",x"49",x"73"),
   502 => (x"70",x"86",x"c4",x"87"),
   503 => (x"87",x"c5",x"05",x"98"),
   504 => (x"e6",x"c0",x"48",x"c0"),
   505 => (x"e6",x"e7",x"c2",x"87"),
   506 => (x"87",x"d2",x"02",x"bf"),
   507 => (x"91",x"c4",x"49",x"74"),
   508 => (x"81",x"de",x"df",x"c2"),
   509 => (x"ff",x"cf",x"4d",x"69"),
   510 => (x"9d",x"ff",x"ff",x"ff"),
   511 => (x"49",x"74",x"87",x"cb"),
   512 => (x"df",x"c2",x"91",x"c2"),
   513 => (x"69",x"9f",x"81",x"de"),
   514 => (x"fe",x"48",x"75",x"4d"),
   515 => (x"5e",x"0e",x"87",x"c6"),
   516 => (x"0e",x"5d",x"5c",x"5b"),
   517 => (x"c0",x"4d",x"71",x"1e"),
   518 => (x"ca",x"49",x"c1",x"1e"),
   519 => (x"86",x"c4",x"87",x"ff"),
   520 => (x"02",x"9c",x"4c",x"70"),
   521 => (x"c2",x"87",x"c0",x"c1"),
   522 => (x"75",x"4a",x"ee",x"e7"),
   523 => (x"87",x"df",x"e0",x"49"),
   524 => (x"c0",x"02",x"98",x"70"),
   525 => (x"4a",x"74",x"87",x"f1"),
   526 => (x"4b",x"cb",x"49",x"75"),
   527 => (x"70",x"87",x"c5",x"e1"),
   528 => (x"e2",x"c0",x"02",x"98"),
   529 => (x"74",x"1e",x"c0",x"87"),
   530 => (x"87",x"c7",x"02",x"9c"),
   531 => (x"c0",x"48",x"a6",x"c4"),
   532 => (x"c4",x"87",x"c5",x"78"),
   533 => (x"78",x"c1",x"48",x"a6"),
   534 => (x"c9",x"49",x"66",x"c4"),
   535 => (x"86",x"c4",x"87",x"ff"),
   536 => (x"05",x"9c",x"4c",x"70"),
   537 => (x"74",x"87",x"c0",x"ff"),
   538 => (x"e7",x"fc",x"26",x"48"),
   539 => (x"5b",x"5e",x"0e",x"87"),
   540 => (x"1e",x"0e",x"5d",x"5c"),
   541 => (x"05",x"9b",x"4b",x"71"),
   542 => (x"48",x"c0",x"87",x"c5"),
   543 => (x"c8",x"87",x"e5",x"c1"),
   544 => (x"7d",x"c0",x"4d",x"a3"),
   545 => (x"c7",x"02",x"66",x"d4"),
   546 => (x"97",x"66",x"d4",x"87"),
   547 => (x"87",x"c5",x"05",x"bf"),
   548 => (x"cf",x"c1",x"48",x"c0"),
   549 => (x"49",x"66",x"d4",x"87"),
   550 => (x"70",x"87",x"f3",x"fd"),
   551 => (x"c1",x"02",x"9c",x"4c"),
   552 => (x"a4",x"dc",x"87",x"c0"),
   553 => (x"da",x"7d",x"69",x"49"),
   554 => (x"a3",x"c4",x"49",x"a4"),
   555 => (x"7a",x"69",x"9f",x"4a"),
   556 => (x"bf",x"e6",x"e7",x"c2"),
   557 => (x"d4",x"87",x"d2",x"02"),
   558 => (x"69",x"9f",x"49",x"a4"),
   559 => (x"ff",x"ff",x"c0",x"49"),
   560 => (x"d0",x"48",x"71",x"99"),
   561 => (x"c2",x"7e",x"70",x"30"),
   562 => (x"6e",x"7e",x"c0",x"87"),
   563 => (x"80",x"6a",x"48",x"49"),
   564 => (x"7b",x"c0",x"7a",x"70"),
   565 => (x"6a",x"49",x"a3",x"cc"),
   566 => (x"49",x"a3",x"d0",x"79"),
   567 => (x"48",x"c1",x"79",x"c0"),
   568 => (x"48",x"c0",x"87",x"c2"),
   569 => (x"87",x"ec",x"fa",x"26"),
   570 => (x"5c",x"5b",x"5e",x"0e"),
   571 => (x"4c",x"71",x"0e",x"5d"),
   572 => (x"ca",x"c1",x"02",x"9c"),
   573 => (x"49",x"a4",x"c8",x"87"),
   574 => (x"c2",x"c1",x"02",x"69"),
   575 => (x"4a",x"66",x"d0",x"87"),
   576 => (x"d4",x"82",x"49",x"6c"),
   577 => (x"66",x"d0",x"5a",x"a6"),
   578 => (x"e7",x"c2",x"b9",x"4d"),
   579 => (x"ff",x"4a",x"bf",x"e2"),
   580 => (x"71",x"99",x"72",x"ba"),
   581 => (x"e4",x"c0",x"02",x"99"),
   582 => (x"4b",x"a4",x"c4",x"87"),
   583 => (x"fb",x"f9",x"49",x"6b"),
   584 => (x"c2",x"7b",x"70",x"87"),
   585 => (x"49",x"bf",x"de",x"e7"),
   586 => (x"7c",x"71",x"81",x"6c"),
   587 => (x"e7",x"c2",x"b9",x"75"),
   588 => (x"ff",x"4a",x"bf",x"e2"),
   589 => (x"71",x"99",x"72",x"ba"),
   590 => (x"dc",x"ff",x"05",x"99"),
   591 => (x"f9",x"7c",x"75",x"87"),
   592 => (x"73",x"1e",x"87",x"d2"),
   593 => (x"9b",x"4b",x"71",x"1e"),
   594 => (x"c8",x"87",x"c7",x"02"),
   595 => (x"05",x"69",x"49",x"a3"),
   596 => (x"48",x"c0",x"87",x"c5"),
   597 => (x"c2",x"87",x"f7",x"c0"),
   598 => (x"4a",x"bf",x"f7",x"eb"),
   599 => (x"69",x"49",x"a3",x"c4"),
   600 => (x"c2",x"89",x"c2",x"49"),
   601 => (x"91",x"bf",x"de",x"e7"),
   602 => (x"c2",x"4a",x"a2",x"71"),
   603 => (x"49",x"bf",x"e2",x"e7"),
   604 => (x"a2",x"71",x"99",x"6b"),
   605 => (x"fc",x"f2",x"c0",x"4a"),
   606 => (x"1e",x"66",x"c8",x"5a"),
   607 => (x"d5",x"ea",x"49",x"72"),
   608 => (x"70",x"86",x"c4",x"87"),
   609 => (x"87",x"c4",x"05",x"98"),
   610 => (x"87",x"c2",x"48",x"c0"),
   611 => (x"c7",x"f8",x"48",x"c1"),
   612 => (x"1e",x"73",x"1e",x"87"),
   613 => (x"02",x"9b",x"4b",x"71"),
   614 => (x"a3",x"c8",x"87",x"c7"),
   615 => (x"c5",x"05",x"69",x"49"),
   616 => (x"c0",x"48",x"c0",x"87"),
   617 => (x"eb",x"c2",x"87",x"f7"),
   618 => (x"c4",x"4a",x"bf",x"f7"),
   619 => (x"49",x"69",x"49",x"a3"),
   620 => (x"e7",x"c2",x"89",x"c2"),
   621 => (x"71",x"91",x"bf",x"de"),
   622 => (x"e7",x"c2",x"4a",x"a2"),
   623 => (x"6b",x"49",x"bf",x"e2"),
   624 => (x"4a",x"a2",x"71",x"99"),
   625 => (x"5a",x"fc",x"f2",x"c0"),
   626 => (x"72",x"1e",x"66",x"c8"),
   627 => (x"87",x"fe",x"e5",x"49"),
   628 => (x"98",x"70",x"86",x"c4"),
   629 => (x"c0",x"87",x"c4",x"05"),
   630 => (x"c1",x"87",x"c2",x"48"),
   631 => (x"87",x"f8",x"f6",x"48"),
   632 => (x"5c",x"5b",x"5e",x"0e"),
   633 => (x"71",x"1e",x"0e",x"5d"),
   634 => (x"4c",x"66",x"d4",x"4b"),
   635 => (x"9b",x"73",x"2c",x"c9"),
   636 => (x"87",x"cf",x"c1",x"02"),
   637 => (x"69",x"49",x"a3",x"c8"),
   638 => (x"87",x"c7",x"c1",x"02"),
   639 => (x"d4",x"4d",x"a3",x"d0"),
   640 => (x"e7",x"c2",x"7d",x"66"),
   641 => (x"ff",x"49",x"bf",x"e2"),
   642 => (x"99",x"4a",x"6b",x"b9"),
   643 => (x"03",x"ac",x"71",x"7e"),
   644 => (x"7b",x"c0",x"87",x"cd"),
   645 => (x"4a",x"a3",x"cc",x"7d"),
   646 => (x"6a",x"49",x"a3",x"c4"),
   647 => (x"72",x"87",x"c2",x"79"),
   648 => (x"02",x"9c",x"74",x"8c"),
   649 => (x"1e",x"49",x"87",x"dd"),
   650 => (x"fb",x"fa",x"49",x"73"),
   651 => (x"d4",x"86",x"c4",x"87"),
   652 => (x"ff",x"c7",x"49",x"66"),
   653 => (x"87",x"cb",x"02",x"99"),
   654 => (x"1e",x"de",x"df",x"c2"),
   655 => (x"c1",x"fc",x"49",x"73"),
   656 => (x"26",x"86",x"c4",x"87"),
   657 => (x"1e",x"87",x"cd",x"f5"),
   658 => (x"4b",x"71",x"1e",x"73"),
   659 => (x"e4",x"c0",x"02",x"9b"),
   660 => (x"cb",x"ec",x"c2",x"87"),
   661 => (x"c2",x"4a",x"73",x"5b"),
   662 => (x"de",x"e7",x"c2",x"8a"),
   663 => (x"c2",x"92",x"49",x"bf"),
   664 => (x"48",x"bf",x"f7",x"eb"),
   665 => (x"ec",x"c2",x"80",x"72"),
   666 => (x"48",x"71",x"58",x"cf"),
   667 => (x"e7",x"c2",x"30",x"c4"),
   668 => (x"ed",x"c0",x"58",x"ee"),
   669 => (x"c7",x"ec",x"c2",x"87"),
   670 => (x"fb",x"eb",x"c2",x"48"),
   671 => (x"ec",x"c2",x"78",x"bf"),
   672 => (x"eb",x"c2",x"48",x"cb"),
   673 => (x"c2",x"78",x"bf",x"ff"),
   674 => (x"02",x"bf",x"e6",x"e7"),
   675 => (x"e7",x"c2",x"87",x"c9"),
   676 => (x"c4",x"49",x"bf",x"de"),
   677 => (x"c2",x"87",x"c7",x"31"),
   678 => (x"49",x"bf",x"c3",x"ec"),
   679 => (x"e7",x"c2",x"31",x"c4"),
   680 => (x"f3",x"f3",x"59",x"ee"),
   681 => (x"5b",x"5e",x"0e",x"87"),
   682 => (x"4a",x"71",x"0e",x"5c"),
   683 => (x"9a",x"72",x"4b",x"c0"),
   684 => (x"87",x"e1",x"c0",x"02"),
   685 => (x"9f",x"49",x"a2",x"da"),
   686 => (x"e7",x"c2",x"4b",x"69"),
   687 => (x"cf",x"02",x"bf",x"e6"),
   688 => (x"49",x"a2",x"d4",x"87"),
   689 => (x"4c",x"49",x"69",x"9f"),
   690 => (x"9c",x"ff",x"ff",x"c0"),
   691 => (x"87",x"c2",x"34",x"d0"),
   692 => (x"49",x"74",x"4c",x"c0"),
   693 => (x"fd",x"49",x"73",x"b3"),
   694 => (x"f9",x"f2",x"87",x"ed"),
   695 => (x"5b",x"5e",x"0e",x"87"),
   696 => (x"f4",x"0e",x"5d",x"5c"),
   697 => (x"c0",x"4a",x"71",x"86"),
   698 => (x"02",x"9a",x"72",x"7e"),
   699 => (x"df",x"c2",x"87",x"d8"),
   700 => (x"78",x"c0",x"48",x"da"),
   701 => (x"48",x"d2",x"df",x"c2"),
   702 => (x"bf",x"cb",x"ec",x"c2"),
   703 => (x"d6",x"df",x"c2",x"78"),
   704 => (x"c7",x"ec",x"c2",x"48"),
   705 => (x"e7",x"c2",x"78",x"bf"),
   706 => (x"50",x"c0",x"48",x"fb"),
   707 => (x"bf",x"ea",x"e7",x"c2"),
   708 => (x"da",x"df",x"c2",x"49"),
   709 => (x"aa",x"71",x"4a",x"bf"),
   710 => (x"87",x"c9",x"c4",x"03"),
   711 => (x"99",x"cf",x"49",x"72"),
   712 => (x"87",x"e9",x"c0",x"05"),
   713 => (x"48",x"f8",x"f2",x"c0"),
   714 => (x"bf",x"d2",x"df",x"c2"),
   715 => (x"de",x"df",x"c2",x"78"),
   716 => (x"d2",x"df",x"c2",x"1e"),
   717 => (x"df",x"c2",x"49",x"bf"),
   718 => (x"a1",x"c1",x"48",x"d2"),
   719 => (x"d5",x"e3",x"71",x"78"),
   720 => (x"c0",x"86",x"c4",x"87"),
   721 => (x"c2",x"48",x"f4",x"f2"),
   722 => (x"cc",x"78",x"de",x"df"),
   723 => (x"f4",x"f2",x"c0",x"87"),
   724 => (x"e0",x"c0",x"48",x"bf"),
   725 => (x"f8",x"f2",x"c0",x"80"),
   726 => (x"da",x"df",x"c2",x"58"),
   727 => (x"80",x"c1",x"48",x"bf"),
   728 => (x"58",x"de",x"df",x"c2"),
   729 => (x"00",x"0c",x"b4",x"27"),
   730 => (x"bf",x"97",x"bf",x"00"),
   731 => (x"c2",x"02",x"9d",x"4d"),
   732 => (x"e5",x"c3",x"87",x"e3"),
   733 => (x"dc",x"c2",x"02",x"ad"),
   734 => (x"f4",x"f2",x"c0",x"87"),
   735 => (x"a3",x"cb",x"4b",x"bf"),
   736 => (x"cf",x"4c",x"11",x"49"),
   737 => (x"d2",x"c1",x"05",x"ac"),
   738 => (x"df",x"49",x"75",x"87"),
   739 => (x"cd",x"89",x"c1",x"99"),
   740 => (x"ee",x"e7",x"c2",x"91"),
   741 => (x"4a",x"a3",x"c1",x"81"),
   742 => (x"a3",x"c3",x"51",x"12"),
   743 => (x"c5",x"51",x"12",x"4a"),
   744 => (x"51",x"12",x"4a",x"a3"),
   745 => (x"12",x"4a",x"a3",x"c7"),
   746 => (x"4a",x"a3",x"c9",x"51"),
   747 => (x"a3",x"ce",x"51",x"12"),
   748 => (x"d0",x"51",x"12",x"4a"),
   749 => (x"51",x"12",x"4a",x"a3"),
   750 => (x"12",x"4a",x"a3",x"d2"),
   751 => (x"4a",x"a3",x"d4",x"51"),
   752 => (x"a3",x"d6",x"51",x"12"),
   753 => (x"d8",x"51",x"12",x"4a"),
   754 => (x"51",x"12",x"4a",x"a3"),
   755 => (x"12",x"4a",x"a3",x"dc"),
   756 => (x"4a",x"a3",x"de",x"51"),
   757 => (x"7e",x"c1",x"51",x"12"),
   758 => (x"74",x"87",x"fa",x"c0"),
   759 => (x"05",x"99",x"c8",x"49"),
   760 => (x"74",x"87",x"eb",x"c0"),
   761 => (x"05",x"99",x"d0",x"49"),
   762 => (x"66",x"dc",x"87",x"d1"),
   763 => (x"87",x"cb",x"c0",x"02"),
   764 => (x"66",x"dc",x"49",x"73"),
   765 => (x"02",x"98",x"70",x"0f"),
   766 => (x"6e",x"87",x"d3",x"c0"),
   767 => (x"87",x"c6",x"c0",x"05"),
   768 => (x"48",x"ee",x"e7",x"c2"),
   769 => (x"f2",x"c0",x"50",x"c0"),
   770 => (x"c2",x"48",x"bf",x"f4"),
   771 => (x"e7",x"c2",x"87",x"e1"),
   772 => (x"50",x"c0",x"48",x"fb"),
   773 => (x"ea",x"e7",x"c2",x"7e"),
   774 => (x"df",x"c2",x"49",x"bf"),
   775 => (x"71",x"4a",x"bf",x"da"),
   776 => (x"f7",x"fb",x"04",x"aa"),
   777 => (x"cb",x"ec",x"c2",x"87"),
   778 => (x"c8",x"c0",x"05",x"bf"),
   779 => (x"e6",x"e7",x"c2",x"87"),
   780 => (x"f8",x"c1",x"02",x"bf"),
   781 => (x"d6",x"df",x"c2",x"87"),
   782 => (x"df",x"ed",x"49",x"bf"),
   783 => (x"c2",x"49",x"70",x"87"),
   784 => (x"c4",x"59",x"da",x"df"),
   785 => (x"df",x"c2",x"48",x"a6"),
   786 => (x"c2",x"78",x"bf",x"d6"),
   787 => (x"02",x"bf",x"e6",x"e7"),
   788 => (x"c4",x"87",x"d8",x"c0"),
   789 => (x"ff",x"cf",x"49",x"66"),
   790 => (x"99",x"f8",x"ff",x"ff"),
   791 => (x"c5",x"c0",x"02",x"a9"),
   792 => (x"c0",x"4c",x"c0",x"87"),
   793 => (x"4c",x"c1",x"87",x"e1"),
   794 => (x"c4",x"87",x"dc",x"c0"),
   795 => (x"ff",x"cf",x"49",x"66"),
   796 => (x"02",x"a9",x"99",x"f8"),
   797 => (x"c8",x"87",x"c8",x"c0"),
   798 => (x"78",x"c0",x"48",x"a6"),
   799 => (x"c8",x"87",x"c5",x"c0"),
   800 => (x"78",x"c1",x"48",x"a6"),
   801 => (x"74",x"4c",x"66",x"c8"),
   802 => (x"e0",x"c0",x"05",x"9c"),
   803 => (x"49",x"66",x"c4",x"87"),
   804 => (x"e7",x"c2",x"89",x"c2"),
   805 => (x"91",x"4a",x"bf",x"de"),
   806 => (x"bf",x"f7",x"eb",x"c2"),
   807 => (x"d2",x"df",x"c2",x"4a"),
   808 => (x"78",x"a1",x"72",x"48"),
   809 => (x"48",x"da",x"df",x"c2"),
   810 => (x"df",x"f9",x"78",x"c0"),
   811 => (x"f4",x"48",x"c0",x"87"),
   812 => (x"87",x"e0",x"eb",x"8e"),
   813 => (x"00",x"00",x"00",x"00"),
   814 => (x"ff",x"ff",x"ff",x"ff"),
   815 => (x"00",x"00",x"0c",x"c4"),
   816 => (x"00",x"00",x"0c",x"cd"),
   817 => (x"33",x"54",x"41",x"46"),
   818 => (x"20",x"20",x"20",x"32"),
   819 => (x"54",x"41",x"46",x"00"),
   820 => (x"20",x"20",x"36",x"31"),
   821 => (x"ff",x"1e",x"00",x"20"),
   822 => (x"ff",x"c3",x"48",x"d4"),
   823 => (x"26",x"48",x"68",x"78"),
   824 => (x"d4",x"ff",x"1e",x"4f"),
   825 => (x"78",x"ff",x"c3",x"48"),
   826 => (x"c0",x"48",x"d0",x"ff"),
   827 => (x"d4",x"ff",x"78",x"e1"),
   828 => (x"c2",x"78",x"d4",x"48"),
   829 => (x"ff",x"48",x"cf",x"ec"),
   830 => (x"26",x"50",x"bf",x"d4"),
   831 => (x"d0",x"ff",x"1e",x"4f"),
   832 => (x"78",x"e0",x"c0",x"48"),
   833 => (x"ff",x"1e",x"4f",x"26"),
   834 => (x"49",x"70",x"87",x"cc"),
   835 => (x"87",x"c6",x"02",x"99"),
   836 => (x"05",x"a9",x"fb",x"c0"),
   837 => (x"48",x"71",x"87",x"f1"),
   838 => (x"5e",x"0e",x"4f",x"26"),
   839 => (x"71",x"0e",x"5c",x"5b"),
   840 => (x"fe",x"4c",x"c0",x"4b"),
   841 => (x"49",x"70",x"87",x"f0"),
   842 => (x"f9",x"c0",x"02",x"99"),
   843 => (x"a9",x"ec",x"c0",x"87"),
   844 => (x"87",x"f2",x"c0",x"02"),
   845 => (x"02",x"a9",x"fb",x"c0"),
   846 => (x"cc",x"87",x"eb",x"c0"),
   847 => (x"03",x"ac",x"b7",x"66"),
   848 => (x"66",x"d0",x"87",x"c7"),
   849 => (x"71",x"87",x"c2",x"02"),
   850 => (x"02",x"99",x"71",x"53"),
   851 => (x"84",x"c1",x"87",x"c2"),
   852 => (x"70",x"87",x"c3",x"fe"),
   853 => (x"cd",x"02",x"99",x"49"),
   854 => (x"a9",x"ec",x"c0",x"87"),
   855 => (x"c0",x"87",x"c7",x"02"),
   856 => (x"ff",x"05",x"a9",x"fb"),
   857 => (x"66",x"d0",x"87",x"d5"),
   858 => (x"c0",x"87",x"c3",x"02"),
   859 => (x"ec",x"c0",x"7b",x"97"),
   860 => (x"87",x"c4",x"05",x"a9"),
   861 => (x"87",x"c5",x"4a",x"74"),
   862 => (x"0a",x"c0",x"4a",x"74"),
   863 => (x"c2",x"48",x"72",x"8a"),
   864 => (x"26",x"4d",x"26",x"87"),
   865 => (x"26",x"4b",x"26",x"4c"),
   866 => (x"c9",x"fd",x"1e",x"4f"),
   867 => (x"c0",x"49",x"70",x"87"),
   868 => (x"04",x"a9",x"b7",x"f0"),
   869 => (x"f9",x"c0",x"87",x"ca"),
   870 => (x"c3",x"01",x"a9",x"b7"),
   871 => (x"89",x"f0",x"c0",x"87"),
   872 => (x"a9",x"b7",x"c1",x"c1"),
   873 => (x"c1",x"87",x"ca",x"04"),
   874 => (x"01",x"a9",x"b7",x"da"),
   875 => (x"f7",x"c0",x"87",x"c3"),
   876 => (x"b7",x"e1",x"c1",x"89"),
   877 => (x"87",x"ca",x"04",x"a9"),
   878 => (x"a9",x"b7",x"fa",x"c1"),
   879 => (x"c0",x"87",x"c3",x"01"),
   880 => (x"48",x"71",x"89",x"fd"),
   881 => (x"5e",x"0e",x"4f",x"26"),
   882 => (x"71",x"0e",x"5c",x"5b"),
   883 => (x"4c",x"d4",x"ff",x"4a"),
   884 => (x"e9",x"c0",x"49",x"72"),
   885 => (x"9b",x"4b",x"70",x"87"),
   886 => (x"c1",x"87",x"c2",x"02"),
   887 => (x"48",x"d0",x"ff",x"8b"),
   888 => (x"d5",x"c1",x"78",x"c5"),
   889 => (x"c6",x"49",x"73",x"7c"),
   890 => (x"fa",x"e2",x"c1",x"31"),
   891 => (x"48",x"4a",x"bf",x"97"),
   892 => (x"7c",x"70",x"b0",x"71"),
   893 => (x"c4",x"48",x"d0",x"ff"),
   894 => (x"fe",x"48",x"73",x"78"),
   895 => (x"5e",x"0e",x"87",x"c5"),
   896 => (x"0e",x"5d",x"5c",x"5b"),
   897 => (x"4c",x"71",x"86",x"f8"),
   898 => (x"d4",x"fb",x"7e",x"c0"),
   899 => (x"c0",x"4b",x"c0",x"87"),
   900 => (x"bf",x"97",x"eb",x"fa"),
   901 => (x"04",x"a9",x"c0",x"49"),
   902 => (x"e9",x"fb",x"87",x"cf"),
   903 => (x"c0",x"83",x"c1",x"87"),
   904 => (x"bf",x"97",x"eb",x"fa"),
   905 => (x"f1",x"06",x"ab",x"49"),
   906 => (x"eb",x"fa",x"c0",x"87"),
   907 => (x"cf",x"02",x"bf",x"97"),
   908 => (x"87",x"e2",x"fa",x"87"),
   909 => (x"02",x"99",x"49",x"70"),
   910 => (x"ec",x"c0",x"87",x"c6"),
   911 => (x"87",x"f1",x"05",x"a9"),
   912 => (x"d1",x"fa",x"4b",x"c0"),
   913 => (x"fa",x"4d",x"70",x"87"),
   914 => (x"a6",x"c8",x"87",x"cc"),
   915 => (x"87",x"c6",x"fa",x"58"),
   916 => (x"83",x"c1",x"4a",x"70"),
   917 => (x"97",x"49",x"a4",x"c8"),
   918 => (x"02",x"ad",x"49",x"69"),
   919 => (x"ff",x"c0",x"87",x"c7"),
   920 => (x"e7",x"c0",x"05",x"ad"),
   921 => (x"49",x"a4",x"c9",x"87"),
   922 => (x"c4",x"49",x"69",x"97"),
   923 => (x"c7",x"02",x"a9",x"66"),
   924 => (x"ff",x"c0",x"48",x"87"),
   925 => (x"87",x"d4",x"05",x"a8"),
   926 => (x"97",x"49",x"a4",x"ca"),
   927 => (x"02",x"aa",x"49",x"69"),
   928 => (x"ff",x"c0",x"87",x"c6"),
   929 => (x"87",x"c4",x"05",x"aa"),
   930 => (x"87",x"d0",x"7e",x"c1"),
   931 => (x"02",x"ad",x"ec",x"c0"),
   932 => (x"fb",x"c0",x"87",x"c6"),
   933 => (x"87",x"c4",x"05",x"ad"),
   934 => (x"7e",x"c1",x"4b",x"c0"),
   935 => (x"e1",x"fe",x"02",x"6e"),
   936 => (x"87",x"d9",x"f9",x"87"),
   937 => (x"8e",x"f8",x"48",x"73"),
   938 => (x"00",x"87",x"d6",x"fb"),
   939 => (x"5c",x"5b",x"5e",x"0e"),
   940 => (x"71",x"1e",x"0e",x"5d"),
   941 => (x"4b",x"d4",x"ff",x"4d"),
   942 => (x"ec",x"c2",x"1e",x"75"),
   943 => (x"ec",x"e6",x"49",x"d4"),
   944 => (x"70",x"86",x"c4",x"87"),
   945 => (x"d5",x"c3",x"02",x"98"),
   946 => (x"dc",x"ec",x"c2",x"87"),
   947 => (x"49",x"75",x"4c",x"bf"),
   948 => (x"ff",x"87",x"f3",x"fb"),
   949 => (x"78",x"c5",x"48",x"d0"),
   950 => (x"c0",x"7b",x"d6",x"c1"),
   951 => (x"49",x"a2",x"75",x"4a"),
   952 => (x"82",x"c1",x"7b",x"11"),
   953 => (x"04",x"aa",x"b7",x"cb"),
   954 => (x"4a",x"cc",x"87",x"f3"),
   955 => (x"c1",x"7b",x"ff",x"c3"),
   956 => (x"b7",x"e0",x"c0",x"82"),
   957 => (x"87",x"f4",x"04",x"aa"),
   958 => (x"c4",x"48",x"d0",x"ff"),
   959 => (x"7b",x"ff",x"c3",x"78"),
   960 => (x"d3",x"c1",x"78",x"c5"),
   961 => (x"c4",x"7b",x"c1",x"7b"),
   962 => (x"02",x"9c",x"74",x"78"),
   963 => (x"c2",x"87",x"ff",x"c1"),
   964 => (x"c8",x"7e",x"de",x"df"),
   965 => (x"c0",x"8c",x"4d",x"c0"),
   966 => (x"c6",x"03",x"ac",x"b7"),
   967 => (x"a4",x"c0",x"c8",x"87"),
   968 => (x"c8",x"4c",x"c0",x"4d"),
   969 => (x"dc",x"05",x"ad",x"c0"),
   970 => (x"cf",x"ec",x"c2",x"87"),
   971 => (x"d0",x"49",x"bf",x"97"),
   972 => (x"87",x"d1",x"02",x"99"),
   973 => (x"ec",x"c2",x"1e",x"c0"),
   974 => (x"c5",x"e8",x"49",x"d4"),
   975 => (x"70",x"86",x"c4",x"87"),
   976 => (x"ee",x"c0",x"4a",x"49"),
   977 => (x"de",x"df",x"c2",x"87"),
   978 => (x"d4",x"ec",x"c2",x"1e"),
   979 => (x"87",x"f2",x"e7",x"49"),
   980 => (x"49",x"70",x"86",x"c4"),
   981 => (x"48",x"d0",x"ff",x"4a"),
   982 => (x"c1",x"78",x"c5",x"c8"),
   983 => (x"97",x"6e",x"7b",x"d4"),
   984 => (x"48",x"6e",x"7b",x"bf"),
   985 => (x"7e",x"70",x"80",x"c1"),
   986 => (x"ff",x"05",x"8d",x"c1"),
   987 => (x"d0",x"ff",x"87",x"f0"),
   988 => (x"72",x"78",x"c4",x"48"),
   989 => (x"87",x"c5",x"05",x"9a"),
   990 => (x"e3",x"c0",x"48",x"c0"),
   991 => (x"c2",x"1e",x"c1",x"87"),
   992 => (x"e5",x"49",x"d4",x"ec"),
   993 => (x"86",x"c4",x"87",x"e2"),
   994 => (x"fe",x"05",x"9c",x"74"),
   995 => (x"d0",x"ff",x"87",x"c1"),
   996 => (x"c1",x"78",x"c5",x"48"),
   997 => (x"7b",x"c0",x"7b",x"d3"),
   998 => (x"48",x"c1",x"78",x"c4"),
   999 => (x"48",x"c0",x"87",x"c2"),
  1000 => (x"26",x"4d",x"26",x"26"),
  1001 => (x"26",x"4b",x"26",x"4c"),
  1002 => (x"5b",x"5e",x"0e",x"4f"),
  1003 => (x"1e",x"0e",x"5d",x"5c"),
  1004 => (x"4c",x"c0",x"4b",x"71"),
  1005 => (x"c0",x"04",x"ab",x"4d"),
  1006 => (x"f7",x"c0",x"87",x"e8"),
  1007 => (x"9d",x"75",x"1e",x"fe"),
  1008 => (x"c0",x"87",x"c4",x"02"),
  1009 => (x"c1",x"87",x"c2",x"4a"),
  1010 => (x"ec",x"49",x"72",x"4a"),
  1011 => (x"86",x"c4",x"87",x"cf"),
  1012 => (x"84",x"c1",x"7e",x"70"),
  1013 => (x"87",x"c2",x"05",x"6e"),
  1014 => (x"85",x"c1",x"4c",x"73"),
  1015 => (x"ff",x"06",x"ac",x"73"),
  1016 => (x"48",x"6e",x"87",x"d8"),
  1017 => (x"87",x"f9",x"fe",x"26"),
  1018 => (x"5c",x"5b",x"5e",x"0e"),
  1019 => (x"cc",x"4b",x"71",x"0e"),
  1020 => (x"87",x"d8",x"02",x"66"),
  1021 => (x"8c",x"f0",x"c0",x"4c"),
  1022 => (x"74",x"87",x"d8",x"02"),
  1023 => (x"02",x"8a",x"c1",x"4a"),
  1024 => (x"02",x"8a",x"87",x"d1"),
  1025 => (x"02",x"8a",x"87",x"cd"),
  1026 => (x"87",x"d9",x"87",x"c9"),
  1027 => (x"db",x"fa",x"49",x"73"),
  1028 => (x"74",x"87",x"d2",x"87"),
  1029 => (x"c1",x"49",x"c0",x"1e"),
  1030 => (x"74",x"87",x"c8",x"db"),
  1031 => (x"c1",x"49",x"73",x"1e"),
  1032 => (x"c8",x"87",x"c0",x"db"),
  1033 => (x"87",x"fb",x"fd",x"86"),
  1034 => (x"5c",x"5b",x"5e",x"0e"),
  1035 => (x"71",x"1e",x"0e",x"5d"),
  1036 => (x"91",x"de",x"49",x"4c"),
  1037 => (x"4d",x"fc",x"ec",x"c2"),
  1038 => (x"6d",x"97",x"85",x"71"),
  1039 => (x"87",x"dc",x"c1",x"02"),
  1040 => (x"bf",x"e8",x"ec",x"c2"),
  1041 => (x"72",x"82",x"74",x"4a"),
  1042 => (x"87",x"dd",x"fd",x"49"),
  1043 => (x"02",x"6e",x"7e",x"70"),
  1044 => (x"c2",x"87",x"f2",x"c0"),
  1045 => (x"6e",x"4b",x"f0",x"ec"),
  1046 => (x"ff",x"49",x"cb",x"4a"),
  1047 => (x"74",x"87",x"c9",x"c1"),
  1048 => (x"c1",x"93",x"cb",x"4b"),
  1049 => (x"c4",x"83",x"ca",x"e3"),
  1050 => (x"e0",x"c2",x"c1",x"83"),
  1051 => (x"c1",x"49",x"74",x"7b"),
  1052 => (x"75",x"87",x"c0",x"c5"),
  1053 => (x"fb",x"e2",x"c1",x"7b"),
  1054 => (x"1e",x"49",x"bf",x"97"),
  1055 => (x"49",x"f0",x"ec",x"c2"),
  1056 => (x"c4",x"87",x"e5",x"fd"),
  1057 => (x"c1",x"49",x"74",x"86"),
  1058 => (x"c0",x"87",x"e8",x"c4"),
  1059 => (x"c7",x"c6",x"c1",x"49"),
  1060 => (x"d0",x"ec",x"c2",x"87"),
  1061 => (x"c1",x"78",x"c0",x"48"),
  1062 => (x"87",x"ff",x"dc",x"49"),
  1063 => (x"87",x"c1",x"fc",x"26"),
  1064 => (x"64",x"61",x"6f",x"4c"),
  1065 => (x"2e",x"67",x"6e",x"69"),
  1066 => (x"0e",x"00",x"2e",x"2e"),
  1067 => (x"0e",x"5c",x"5b",x"5e"),
  1068 => (x"c2",x"4a",x"4b",x"71"),
  1069 => (x"82",x"bf",x"e8",x"ec"),
  1070 => (x"ec",x"fb",x"49",x"72"),
  1071 => (x"9c",x"4c",x"70",x"87"),
  1072 => (x"49",x"87",x"c4",x"02"),
  1073 => (x"c2",x"87",x"de",x"e7"),
  1074 => (x"c0",x"48",x"e8",x"ec"),
  1075 => (x"dc",x"49",x"c1",x"78"),
  1076 => (x"ce",x"fb",x"87",x"c9"),
  1077 => (x"5b",x"5e",x"0e",x"87"),
  1078 => (x"f4",x"0e",x"5d",x"5c"),
  1079 => (x"de",x"df",x"c2",x"86"),
  1080 => (x"c4",x"4c",x"c0",x"4d"),
  1081 => (x"78",x"c0",x"48",x"a6"),
  1082 => (x"bf",x"e8",x"ec",x"c2"),
  1083 => (x"06",x"a9",x"c0",x"49"),
  1084 => (x"c2",x"87",x"c1",x"c1"),
  1085 => (x"98",x"48",x"de",x"df"),
  1086 => (x"87",x"f8",x"c0",x"02"),
  1087 => (x"1e",x"fe",x"f7",x"c0"),
  1088 => (x"c7",x"02",x"66",x"c8"),
  1089 => (x"48",x"a6",x"c4",x"87"),
  1090 => (x"87",x"c5",x"78",x"c0"),
  1091 => (x"c1",x"48",x"a6",x"c4"),
  1092 => (x"49",x"66",x"c4",x"78"),
  1093 => (x"c4",x"87",x"c6",x"e7"),
  1094 => (x"c1",x"4d",x"70",x"86"),
  1095 => (x"48",x"66",x"c4",x"84"),
  1096 => (x"a6",x"c8",x"80",x"c1"),
  1097 => (x"e8",x"ec",x"c2",x"58"),
  1098 => (x"03",x"ac",x"49",x"bf"),
  1099 => (x"9d",x"75",x"87",x"c6"),
  1100 => (x"87",x"c8",x"ff",x"05"),
  1101 => (x"9d",x"75",x"4c",x"c0"),
  1102 => (x"87",x"e0",x"c3",x"02"),
  1103 => (x"1e",x"fe",x"f7",x"c0"),
  1104 => (x"c7",x"02",x"66",x"c8"),
  1105 => (x"48",x"a6",x"cc",x"87"),
  1106 => (x"87",x"c5",x"78",x"c0"),
  1107 => (x"c1",x"48",x"a6",x"cc"),
  1108 => (x"49",x"66",x"cc",x"78"),
  1109 => (x"c4",x"87",x"c6",x"e6"),
  1110 => (x"6e",x"7e",x"70",x"86"),
  1111 => (x"87",x"e9",x"c2",x"02"),
  1112 => (x"81",x"cb",x"49",x"6e"),
  1113 => (x"d0",x"49",x"69",x"97"),
  1114 => (x"d6",x"c1",x"02",x"99"),
  1115 => (x"eb",x"c2",x"c1",x"87"),
  1116 => (x"cb",x"49",x"74",x"4a"),
  1117 => (x"ca",x"e3",x"c1",x"91"),
  1118 => (x"c8",x"79",x"72",x"81"),
  1119 => (x"51",x"ff",x"c3",x"81"),
  1120 => (x"91",x"de",x"49",x"74"),
  1121 => (x"4d",x"fc",x"ec",x"c2"),
  1122 => (x"c1",x"c2",x"85",x"71"),
  1123 => (x"a5",x"c1",x"7d",x"97"),
  1124 => (x"51",x"e0",x"c0",x"49"),
  1125 => (x"97",x"ee",x"e7",x"c2"),
  1126 => (x"87",x"d2",x"02",x"bf"),
  1127 => (x"a5",x"c2",x"84",x"c1"),
  1128 => (x"ee",x"e7",x"c2",x"4b"),
  1129 => (x"fe",x"49",x"db",x"4a"),
  1130 => (x"c1",x"87",x"fd",x"fb"),
  1131 => (x"a5",x"cd",x"87",x"db"),
  1132 => (x"c1",x"51",x"c0",x"49"),
  1133 => (x"4b",x"a5",x"c2",x"84"),
  1134 => (x"49",x"cb",x"4a",x"6e"),
  1135 => (x"87",x"e8",x"fb",x"fe"),
  1136 => (x"c1",x"87",x"c6",x"c1"),
  1137 => (x"74",x"4a",x"e8",x"c0"),
  1138 => (x"c1",x"91",x"cb",x"49"),
  1139 => (x"72",x"81",x"ca",x"e3"),
  1140 => (x"ee",x"e7",x"c2",x"79"),
  1141 => (x"d8",x"02",x"bf",x"97"),
  1142 => (x"de",x"49",x"74",x"87"),
  1143 => (x"c2",x"84",x"c1",x"91"),
  1144 => (x"71",x"4b",x"fc",x"ec"),
  1145 => (x"ee",x"e7",x"c2",x"83"),
  1146 => (x"fe",x"49",x"dd",x"4a"),
  1147 => (x"d8",x"87",x"f9",x"fa"),
  1148 => (x"de",x"4b",x"74",x"87"),
  1149 => (x"fc",x"ec",x"c2",x"93"),
  1150 => (x"49",x"a3",x"cb",x"83"),
  1151 => (x"84",x"c1",x"51",x"c0"),
  1152 => (x"cb",x"4a",x"6e",x"73"),
  1153 => (x"df",x"fa",x"fe",x"49"),
  1154 => (x"48",x"66",x"c4",x"87"),
  1155 => (x"a6",x"c8",x"80",x"c1"),
  1156 => (x"03",x"ac",x"c7",x"58"),
  1157 => (x"6e",x"87",x"c5",x"c0"),
  1158 => (x"87",x"e0",x"fc",x"05"),
  1159 => (x"8e",x"f4",x"48",x"74"),
  1160 => (x"1e",x"87",x"fe",x"f5"),
  1161 => (x"4b",x"71",x"1e",x"73"),
  1162 => (x"c1",x"91",x"cb",x"49"),
  1163 => (x"c8",x"81",x"ca",x"e3"),
  1164 => (x"e2",x"c1",x"4a",x"a1"),
  1165 => (x"50",x"12",x"48",x"fa"),
  1166 => (x"c0",x"4a",x"a1",x"c9"),
  1167 => (x"12",x"48",x"eb",x"fa"),
  1168 => (x"c1",x"81",x"ca",x"50"),
  1169 => (x"11",x"48",x"fb",x"e2"),
  1170 => (x"fb",x"e2",x"c1",x"50"),
  1171 => (x"1e",x"49",x"bf",x"97"),
  1172 => (x"d3",x"f6",x"49",x"c0"),
  1173 => (x"d0",x"ec",x"c2",x"87"),
  1174 => (x"c1",x"78",x"de",x"48"),
  1175 => (x"87",x"fb",x"d5",x"49"),
  1176 => (x"87",x"c1",x"f5",x"26"),
  1177 => (x"49",x"4a",x"71",x"1e"),
  1178 => (x"e3",x"c1",x"91",x"cb"),
  1179 => (x"81",x"c8",x"81",x"ca"),
  1180 => (x"ec",x"c2",x"48",x"11"),
  1181 => (x"ec",x"c2",x"58",x"d4"),
  1182 => (x"78",x"c0",x"48",x"e8"),
  1183 => (x"da",x"d5",x"49",x"c1"),
  1184 => (x"1e",x"4f",x"26",x"87"),
  1185 => (x"fe",x"c0",x"49",x"c0"),
  1186 => (x"4f",x"26",x"87",x"ce"),
  1187 => (x"02",x"99",x"71",x"1e"),
  1188 => (x"e4",x"c1",x"87",x"d2"),
  1189 => (x"50",x"c0",x"48",x"df"),
  1190 => (x"c9",x"c1",x"80",x"f7"),
  1191 => (x"e3",x"c1",x"40",x"e4"),
  1192 => (x"87",x"ce",x"78",x"c3"),
  1193 => (x"48",x"db",x"e4",x"c1"),
  1194 => (x"78",x"fc",x"e2",x"c1"),
  1195 => (x"ca",x"c1",x"80",x"fc"),
  1196 => (x"4f",x"26",x"78",x"c3"),
  1197 => (x"5c",x"5b",x"5e",x"0e"),
  1198 => (x"4a",x"4c",x"71",x"0e"),
  1199 => (x"e3",x"c1",x"92",x"cb"),
  1200 => (x"a2",x"c8",x"82",x"ca"),
  1201 => (x"4b",x"a2",x"c9",x"49"),
  1202 => (x"1e",x"4b",x"6b",x"97"),
  1203 => (x"1e",x"49",x"69",x"97"),
  1204 => (x"49",x"12",x"82",x"ca"),
  1205 => (x"87",x"c7",x"e7",x"c0"),
  1206 => (x"fe",x"d3",x"49",x"c0"),
  1207 => (x"c0",x"49",x"74",x"87"),
  1208 => (x"f8",x"87",x"d0",x"fb"),
  1209 => (x"87",x"fb",x"f2",x"8e"),
  1210 => (x"71",x"1e",x"73",x"1e"),
  1211 => (x"c3",x"ff",x"49",x"4b"),
  1212 => (x"fe",x"49",x"73",x"87"),
  1213 => (x"ec",x"f2",x"87",x"fe"),
  1214 => (x"1e",x"73",x"1e",x"87"),
  1215 => (x"a3",x"c6",x"4b",x"71"),
  1216 => (x"87",x"db",x"02",x"4a"),
  1217 => (x"d6",x"02",x"8a",x"c1"),
  1218 => (x"c1",x"02",x"8a",x"87"),
  1219 => (x"02",x"8a",x"87",x"da"),
  1220 => (x"8a",x"87",x"fc",x"c0"),
  1221 => (x"87",x"e1",x"c0",x"02"),
  1222 => (x"87",x"cb",x"02",x"8a"),
  1223 => (x"c7",x"87",x"db",x"c1"),
  1224 => (x"87",x"c0",x"fd",x"49"),
  1225 => (x"c2",x"87",x"de",x"c1"),
  1226 => (x"02",x"bf",x"e8",x"ec"),
  1227 => (x"48",x"87",x"cb",x"c1"),
  1228 => (x"ec",x"c2",x"88",x"c1"),
  1229 => (x"c1",x"c1",x"58",x"ec"),
  1230 => (x"ec",x"ec",x"c2",x"87"),
  1231 => (x"f9",x"c0",x"02",x"bf"),
  1232 => (x"e8",x"ec",x"c2",x"87"),
  1233 => (x"80",x"c1",x"48",x"bf"),
  1234 => (x"58",x"ec",x"ec",x"c2"),
  1235 => (x"c2",x"87",x"eb",x"c0"),
  1236 => (x"49",x"bf",x"e8",x"ec"),
  1237 => (x"ec",x"c2",x"89",x"c6"),
  1238 => (x"b7",x"c0",x"59",x"ec"),
  1239 => (x"87",x"da",x"03",x"a9"),
  1240 => (x"48",x"e8",x"ec",x"c2"),
  1241 => (x"87",x"d2",x"78",x"c0"),
  1242 => (x"bf",x"ec",x"ec",x"c2"),
  1243 => (x"c2",x"87",x"cb",x"02"),
  1244 => (x"48",x"bf",x"e8",x"ec"),
  1245 => (x"ec",x"c2",x"80",x"c6"),
  1246 => (x"49",x"c0",x"58",x"ec"),
  1247 => (x"73",x"87",x"dc",x"d1"),
  1248 => (x"ee",x"f8",x"c0",x"49"),
  1249 => (x"87",x"dd",x"f0",x"87"),
  1250 => (x"5c",x"5b",x"5e",x"0e"),
  1251 => (x"cc",x"4c",x"71",x"0e"),
  1252 => (x"4b",x"74",x"1e",x"66"),
  1253 => (x"e3",x"c1",x"93",x"cb"),
  1254 => (x"a3",x"c4",x"83",x"ca"),
  1255 => (x"fe",x"49",x"6a",x"4a"),
  1256 => (x"c1",x"87",x"d5",x"f4"),
  1257 => (x"c8",x"7b",x"e3",x"c8"),
  1258 => (x"66",x"d4",x"49",x"a3"),
  1259 => (x"49",x"a3",x"c9",x"51"),
  1260 => (x"ca",x"51",x"66",x"d8"),
  1261 => (x"66",x"dc",x"49",x"a3"),
  1262 => (x"e6",x"ef",x"26",x"51"),
  1263 => (x"5b",x"5e",x"0e",x"87"),
  1264 => (x"ff",x"0e",x"5d",x"5c"),
  1265 => (x"a6",x"d8",x"86",x"d0"),
  1266 => (x"48",x"a6",x"c4",x"59"),
  1267 => (x"80",x"c4",x"78",x"c0"),
  1268 => (x"78",x"66",x"c4",x"c1"),
  1269 => (x"78",x"c1",x"80",x"c4"),
  1270 => (x"78",x"c1",x"80",x"c4"),
  1271 => (x"48",x"ec",x"ec",x"c2"),
  1272 => (x"ec",x"c2",x"78",x"c1"),
  1273 => (x"de",x"48",x"bf",x"d0"),
  1274 => (x"87",x"cb",x"05",x"a8"),
  1275 => (x"70",x"87",x"e6",x"f3"),
  1276 => (x"59",x"a6",x"c8",x"49"),
  1277 => (x"e3",x"87",x"ec",x"ce"),
  1278 => (x"c9",x"e4",x"87",x"e7"),
  1279 => (x"87",x"d6",x"e3",x"87"),
  1280 => (x"fb",x"c0",x"4c",x"70"),
  1281 => (x"d0",x"c1",x"02",x"ac"),
  1282 => (x"05",x"66",x"d4",x"87"),
  1283 => (x"c0",x"87",x"c2",x"c1"),
  1284 => (x"1e",x"c1",x"1e",x"1e"),
  1285 => (x"1e",x"fd",x"e4",x"c1"),
  1286 => (x"eb",x"fd",x"49",x"c0"),
  1287 => (x"66",x"d0",x"c1",x"87"),
  1288 => (x"6a",x"82",x"c4",x"4a"),
  1289 => (x"74",x"81",x"c7",x"49"),
  1290 => (x"d8",x"1e",x"c1",x"51"),
  1291 => (x"c8",x"49",x"6a",x"1e"),
  1292 => (x"87",x"e6",x"e3",x"81"),
  1293 => (x"c4",x"c1",x"86",x"d8"),
  1294 => (x"a8",x"c0",x"48",x"66"),
  1295 => (x"c4",x"87",x"c7",x"01"),
  1296 => (x"78",x"c1",x"48",x"a6"),
  1297 => (x"c4",x"c1",x"87",x"ce"),
  1298 => (x"88",x"c1",x"48",x"66"),
  1299 => (x"c3",x"58",x"a6",x"cc"),
  1300 => (x"87",x"f2",x"e2",x"87"),
  1301 => (x"c2",x"48",x"a6",x"cc"),
  1302 => (x"02",x"9c",x"74",x"78"),
  1303 => (x"c4",x"87",x"c0",x"cd"),
  1304 => (x"c8",x"c1",x"48",x"66"),
  1305 => (x"cc",x"03",x"a8",x"66"),
  1306 => (x"a6",x"d8",x"87",x"f5"),
  1307 => (x"c4",x"78",x"c0",x"48"),
  1308 => (x"e1",x"78",x"c0",x"80"),
  1309 => (x"4c",x"70",x"87",x"e0"),
  1310 => (x"05",x"ac",x"d0",x"c1"),
  1311 => (x"dc",x"87",x"d8",x"c2"),
  1312 => (x"c4",x"e4",x"7e",x"66"),
  1313 => (x"c0",x"49",x"70",x"87"),
  1314 => (x"e1",x"59",x"a6",x"e0"),
  1315 => (x"4c",x"70",x"87",x"c8"),
  1316 => (x"05",x"ac",x"ec",x"c0"),
  1317 => (x"c4",x"87",x"eb",x"c1"),
  1318 => (x"91",x"cb",x"49",x"66"),
  1319 => (x"81",x"66",x"c0",x"c1"),
  1320 => (x"6a",x"4a",x"a1",x"c4"),
  1321 => (x"4a",x"a1",x"c8",x"4d"),
  1322 => (x"c1",x"52",x"66",x"dc"),
  1323 => (x"e0",x"79",x"e4",x"c9"),
  1324 => (x"4c",x"70",x"87",x"e4"),
  1325 => (x"87",x"d8",x"02",x"9c"),
  1326 => (x"02",x"ac",x"fb",x"c0"),
  1327 => (x"55",x"74",x"87",x"d2"),
  1328 => (x"70",x"87",x"d3",x"e0"),
  1329 => (x"c7",x"02",x"9c",x"4c"),
  1330 => (x"ac",x"fb",x"c0",x"87"),
  1331 => (x"87",x"ee",x"ff",x"05"),
  1332 => (x"c2",x"55",x"e0",x"c0"),
  1333 => (x"97",x"c0",x"55",x"c1"),
  1334 => (x"49",x"66",x"d4",x"7d"),
  1335 => (x"db",x"05",x"a9",x"6e"),
  1336 => (x"48",x"66",x"c4",x"87"),
  1337 => (x"04",x"a8",x"66",x"c8"),
  1338 => (x"66",x"c4",x"87",x"ca"),
  1339 => (x"c8",x"80",x"c1",x"48"),
  1340 => (x"87",x"c8",x"58",x"a6"),
  1341 => (x"c1",x"48",x"66",x"c8"),
  1342 => (x"58",x"a6",x"cc",x"88"),
  1343 => (x"87",x"d6",x"df",x"ff"),
  1344 => (x"d0",x"c1",x"4c",x"70"),
  1345 => (x"87",x"c8",x"05",x"ac"),
  1346 => (x"c1",x"48",x"66",x"d0"),
  1347 => (x"58",x"a6",x"d4",x"80"),
  1348 => (x"02",x"ac",x"d0",x"c1"),
  1349 => (x"c0",x"87",x"e8",x"fd"),
  1350 => (x"d4",x"48",x"a6",x"e0"),
  1351 => (x"66",x"dc",x"78",x"66"),
  1352 => (x"66",x"e0",x"c0",x"48"),
  1353 => (x"c8",x"c9",x"05",x"a8"),
  1354 => (x"a6",x"e4",x"c0",x"87"),
  1355 => (x"7e",x"78",x"c0",x"48"),
  1356 => (x"fb",x"c0",x"48",x"74"),
  1357 => (x"a6",x"ec",x"c0",x"88"),
  1358 => (x"02",x"98",x"70",x"58"),
  1359 => (x"48",x"87",x"cd",x"c8"),
  1360 => (x"ec",x"c0",x"88",x"cb"),
  1361 => (x"98",x"70",x"58",x"a6"),
  1362 => (x"87",x"d2",x"c1",x"02"),
  1363 => (x"c0",x"88",x"c9",x"48"),
  1364 => (x"70",x"58",x"a6",x"ec"),
  1365 => (x"db",x"c3",x"02",x"98"),
  1366 => (x"88",x"c4",x"48",x"87"),
  1367 => (x"58",x"a6",x"ec",x"c0"),
  1368 => (x"d0",x"02",x"98",x"70"),
  1369 => (x"88",x"c1",x"48",x"87"),
  1370 => (x"58",x"a6",x"ec",x"c0"),
  1371 => (x"c3",x"02",x"98",x"70"),
  1372 => (x"d1",x"c7",x"87",x"c2"),
  1373 => (x"48",x"a6",x"d8",x"87"),
  1374 => (x"ff",x"78",x"f0",x"c0"),
  1375 => (x"70",x"87",x"d7",x"dd"),
  1376 => (x"ac",x"ec",x"c0",x"4c"),
  1377 => (x"87",x"c3",x"c0",x"02"),
  1378 => (x"c0",x"5c",x"a6",x"dc"),
  1379 => (x"cd",x"02",x"ac",x"ec"),
  1380 => (x"c1",x"dd",x"ff",x"87"),
  1381 => (x"c0",x"4c",x"70",x"87"),
  1382 => (x"ff",x"05",x"ac",x"ec"),
  1383 => (x"ec",x"c0",x"87",x"f3"),
  1384 => (x"c4",x"c0",x"02",x"ac"),
  1385 => (x"ed",x"dc",x"ff",x"87"),
  1386 => (x"1e",x"66",x"d8",x"87"),
  1387 => (x"1e",x"49",x"66",x"d4"),
  1388 => (x"1e",x"49",x"66",x"d4"),
  1389 => (x"1e",x"fd",x"e4",x"c1"),
  1390 => (x"f7",x"49",x"66",x"d4"),
  1391 => (x"1e",x"c0",x"87",x"ca"),
  1392 => (x"66",x"dc",x"1e",x"ca"),
  1393 => (x"c1",x"91",x"cb",x"49"),
  1394 => (x"d8",x"81",x"66",x"d8"),
  1395 => (x"a1",x"c4",x"48",x"a6"),
  1396 => (x"bf",x"66",x"d8",x"78"),
  1397 => (x"c1",x"dd",x"ff",x"49"),
  1398 => (x"c0",x"86",x"d8",x"87"),
  1399 => (x"c1",x"06",x"a8",x"b7"),
  1400 => (x"1e",x"c1",x"87",x"c5"),
  1401 => (x"66",x"c8",x"1e",x"de"),
  1402 => (x"dc",x"ff",x"49",x"bf"),
  1403 => (x"86",x"c8",x"87",x"ec"),
  1404 => (x"c0",x"48",x"49",x"70"),
  1405 => (x"a6",x"dc",x"88",x"08"),
  1406 => (x"a8",x"b7",x"c0",x"58"),
  1407 => (x"87",x"e7",x"c0",x"06"),
  1408 => (x"dd",x"48",x"66",x"d8"),
  1409 => (x"de",x"03",x"a8",x"b7"),
  1410 => (x"49",x"bf",x"6e",x"87"),
  1411 => (x"c0",x"81",x"66",x"d8"),
  1412 => (x"66",x"d8",x"51",x"e0"),
  1413 => (x"6e",x"81",x"c1",x"49"),
  1414 => (x"c1",x"c2",x"81",x"bf"),
  1415 => (x"49",x"66",x"d8",x"51"),
  1416 => (x"bf",x"6e",x"81",x"c2"),
  1417 => (x"cc",x"51",x"c0",x"81"),
  1418 => (x"80",x"c1",x"48",x"66"),
  1419 => (x"c1",x"58",x"a6",x"d0"),
  1420 => (x"87",x"d8",x"c4",x"7e"),
  1421 => (x"87",x"d1",x"dd",x"ff"),
  1422 => (x"ff",x"58",x"a6",x"dc"),
  1423 => (x"c0",x"87",x"ca",x"dd"),
  1424 => (x"c0",x"58",x"a6",x"ec"),
  1425 => (x"c0",x"05",x"a8",x"ec"),
  1426 => (x"e8",x"c0",x"87",x"ca"),
  1427 => (x"66",x"d8",x"48",x"a6"),
  1428 => (x"87",x"c4",x"c0",x"78"),
  1429 => (x"87",x"fe",x"d9",x"ff"),
  1430 => (x"cb",x"49",x"66",x"c4"),
  1431 => (x"66",x"c0",x"c1",x"91"),
  1432 => (x"70",x"80",x"71",x"48"),
  1433 => (x"c8",x"49",x"6e",x"7e"),
  1434 => (x"ca",x"4a",x"6e",x"81"),
  1435 => (x"52",x"66",x"d8",x"82"),
  1436 => (x"4a",x"66",x"e8",x"c0"),
  1437 => (x"66",x"d8",x"82",x"c1"),
  1438 => (x"72",x"48",x"c1",x"8a"),
  1439 => (x"c1",x"4a",x"70",x"30"),
  1440 => (x"79",x"97",x"72",x"8a"),
  1441 => (x"1e",x"49",x"69",x"97"),
  1442 => (x"d7",x"49",x"66",x"dc"),
  1443 => (x"86",x"c4",x"87",x"d3"),
  1444 => (x"58",x"a6",x"f0",x"c0"),
  1445 => (x"81",x"c4",x"49",x"6e"),
  1446 => (x"e0",x"c0",x"4d",x"69"),
  1447 => (x"66",x"dc",x"48",x"66"),
  1448 => (x"c8",x"c0",x"02",x"a8"),
  1449 => (x"48",x"a6",x"d8",x"87"),
  1450 => (x"c5",x"c0",x"78",x"c0"),
  1451 => (x"48",x"a6",x"d8",x"87"),
  1452 => (x"66",x"d8",x"78",x"c1"),
  1453 => (x"1e",x"e0",x"c0",x"1e"),
  1454 => (x"d9",x"ff",x"49",x"75"),
  1455 => (x"86",x"c8",x"87",x"dc"),
  1456 => (x"b7",x"c0",x"4c",x"70"),
  1457 => (x"d4",x"c1",x"06",x"ac"),
  1458 => (x"c0",x"85",x"74",x"87"),
  1459 => (x"89",x"74",x"49",x"e0"),
  1460 => (x"df",x"c1",x"4b",x"75"),
  1461 => (x"fe",x"71",x"4a",x"d8"),
  1462 => (x"c2",x"87",x"cd",x"e7"),
  1463 => (x"66",x"e4",x"c0",x"85"),
  1464 => (x"c0",x"80",x"c1",x"48"),
  1465 => (x"c0",x"58",x"a6",x"e8"),
  1466 => (x"c1",x"49",x"66",x"ec"),
  1467 => (x"02",x"a9",x"70",x"81"),
  1468 => (x"d8",x"87",x"c8",x"c0"),
  1469 => (x"78",x"c0",x"48",x"a6"),
  1470 => (x"d8",x"87",x"c5",x"c0"),
  1471 => (x"78",x"c1",x"48",x"a6"),
  1472 => (x"c2",x"1e",x"66",x"d8"),
  1473 => (x"e0",x"c0",x"49",x"a4"),
  1474 => (x"70",x"88",x"71",x"48"),
  1475 => (x"49",x"75",x"1e",x"49"),
  1476 => (x"87",x"c6",x"d8",x"ff"),
  1477 => (x"b7",x"c0",x"86",x"c8"),
  1478 => (x"c0",x"ff",x"01",x"a8"),
  1479 => (x"66",x"e4",x"c0",x"87"),
  1480 => (x"87",x"d1",x"c0",x"02"),
  1481 => (x"81",x"c9",x"49",x"6e"),
  1482 => (x"51",x"66",x"e4",x"c0"),
  1483 => (x"ca",x"c1",x"48",x"6e"),
  1484 => (x"cc",x"c0",x"78",x"f4"),
  1485 => (x"c9",x"49",x"6e",x"87"),
  1486 => (x"6e",x"51",x"c2",x"81"),
  1487 => (x"e8",x"cb",x"c1",x"48"),
  1488 => (x"c0",x"7e",x"c1",x"78"),
  1489 => (x"d6",x"ff",x"87",x"c6"),
  1490 => (x"4c",x"70",x"87",x"fc"),
  1491 => (x"f5",x"c0",x"02",x"6e"),
  1492 => (x"48",x"66",x"c4",x"87"),
  1493 => (x"04",x"a8",x"66",x"c8"),
  1494 => (x"c4",x"87",x"cb",x"c0"),
  1495 => (x"80",x"c1",x"48",x"66"),
  1496 => (x"c0",x"58",x"a6",x"c8"),
  1497 => (x"66",x"c8",x"87",x"e0"),
  1498 => (x"cc",x"88",x"c1",x"48"),
  1499 => (x"d5",x"c0",x"58",x"a6"),
  1500 => (x"ac",x"c6",x"c1",x"87"),
  1501 => (x"87",x"c8",x"c0",x"05"),
  1502 => (x"c1",x"48",x"66",x"cc"),
  1503 => (x"58",x"a6",x"d0",x"80"),
  1504 => (x"87",x"c2",x"d6",x"ff"),
  1505 => (x"66",x"d0",x"4c",x"70"),
  1506 => (x"d4",x"80",x"c1",x"48"),
  1507 => (x"9c",x"74",x"58",x"a6"),
  1508 => (x"87",x"cb",x"c0",x"02"),
  1509 => (x"c1",x"48",x"66",x"c4"),
  1510 => (x"04",x"a8",x"66",x"c8"),
  1511 => (x"ff",x"87",x"cb",x"f3"),
  1512 => (x"c4",x"87",x"da",x"d5"),
  1513 => (x"a8",x"c7",x"48",x"66"),
  1514 => (x"87",x"e5",x"c0",x"03"),
  1515 => (x"48",x"ec",x"ec",x"c2"),
  1516 => (x"66",x"c4",x"78",x"c0"),
  1517 => (x"c1",x"91",x"cb",x"49"),
  1518 => (x"c4",x"81",x"66",x"c0"),
  1519 => (x"4a",x"6a",x"4a",x"a1"),
  1520 => (x"c4",x"79",x"52",x"c0"),
  1521 => (x"80",x"c1",x"48",x"66"),
  1522 => (x"c7",x"58",x"a6",x"c8"),
  1523 => (x"db",x"ff",x"04",x"a8"),
  1524 => (x"8e",x"d0",x"ff",x"87"),
  1525 => (x"87",x"c9",x"df",x"ff"),
  1526 => (x"1e",x"00",x"20",x"3a"),
  1527 => (x"4b",x"71",x"1e",x"73"),
  1528 => (x"87",x"c6",x"02",x"9b"),
  1529 => (x"48",x"e8",x"ec",x"c2"),
  1530 => (x"1e",x"c7",x"78",x"c0"),
  1531 => (x"bf",x"e8",x"ec",x"c2"),
  1532 => (x"e3",x"c1",x"1e",x"49"),
  1533 => (x"ec",x"c2",x"1e",x"ca"),
  1534 => (x"ee",x"49",x"bf",x"d0"),
  1535 => (x"86",x"cc",x"87",x"ff"),
  1536 => (x"bf",x"d0",x"ec",x"c2"),
  1537 => (x"87",x"c4",x"ea",x"49"),
  1538 => (x"c8",x"02",x"9b",x"73"),
  1539 => (x"ca",x"e3",x"c1",x"87"),
  1540 => (x"f0",x"e7",x"c0",x"49"),
  1541 => (x"cc",x"de",x"ff",x"87"),
  1542 => (x"e2",x"c1",x"1e",x"87"),
  1543 => (x"50",x"c0",x"48",x"fa"),
  1544 => (x"bf",x"ed",x"e4",x"c1"),
  1545 => (x"c3",x"da",x"ff",x"49"),
  1546 => (x"26",x"48",x"c0",x"87"),
  1547 => (x"eb",x"c7",x"1e",x"4f"),
  1548 => (x"fe",x"49",x"c1",x"87"),
  1549 => (x"ea",x"fe",x"87",x"e5"),
  1550 => (x"98",x"70",x"87",x"e3"),
  1551 => (x"fe",x"87",x"cd",x"02"),
  1552 => (x"70",x"87",x"de",x"f3"),
  1553 => (x"87",x"c4",x"02",x"98"),
  1554 => (x"87",x"c2",x"4a",x"c1"),
  1555 => (x"9a",x"72",x"4a",x"c0"),
  1556 => (x"c0",x"87",x"ce",x"05"),
  1557 => (x"c1",x"e2",x"c1",x"1e"),
  1558 => (x"c0",x"f3",x"c0",x"49"),
  1559 => (x"fe",x"86",x"c4",x"87"),
  1560 => (x"e8",x"fc",x"c0",x"87"),
  1561 => (x"c1",x"1e",x"c0",x"87"),
  1562 => (x"c0",x"49",x"cc",x"e2"),
  1563 => (x"c0",x"87",x"ee",x"f2"),
  1564 => (x"87",x"e5",x"fe",x"1e"),
  1565 => (x"f2",x"c0",x"49",x"70"),
  1566 => (x"de",x"c3",x"87",x"e3"),
  1567 => (x"26",x"8e",x"f8",x"87"),
  1568 => (x"20",x"44",x"53",x"4f"),
  1569 => (x"6c",x"69",x"61",x"66"),
  1570 => (x"00",x"2e",x"64",x"65"),
  1571 => (x"74",x"6f",x"6f",x"42"),
  1572 => (x"2e",x"67",x"6e",x"69"),
  1573 => (x"1e",x"00",x"2e",x"2e"),
  1574 => (x"87",x"c5",x"ea",x"c0"),
  1575 => (x"87",x"f3",x"f5",x"c0"),
  1576 => (x"4f",x"26",x"87",x"f6"),
  1577 => (x"e8",x"ec",x"c2",x"1e"),
  1578 => (x"c2",x"78",x"c0",x"48"),
  1579 => (x"c0",x"48",x"d0",x"ec"),
  1580 => (x"87",x"f9",x"fd",x"78"),
  1581 => (x"48",x"c0",x"87",x"e1"),
  1582 => (x"00",x"00",x"4f",x"26"),
  1583 => (x"78",x"45",x"20",x"80"),
  1584 => (x"80",x"00",x"74",x"69"),
  1585 => (x"63",x"61",x"42",x"20"),
  1586 => (x"12",x"64",x"00",x"6b"),
  1587 => (x"2b",x"3c",x"00",x"00"),
  1588 => (x"00",x"00",x"00",x"00"),
  1589 => (x"00",x"12",x"64",x"00"),
  1590 => (x"00",x"2b",x"5a",x"00"),
  1591 => (x"00",x"00",x"00",x"00"),
  1592 => (x"00",x"00",x"12",x"64"),
  1593 => (x"00",x"00",x"2b",x"78"),
  1594 => (x"64",x"00",x"00",x"00"),
  1595 => (x"96",x"00",x"00",x"12"),
  1596 => (x"00",x"00",x"00",x"2b"),
  1597 => (x"12",x"64",x"00",x"00"),
  1598 => (x"2b",x"b4",x"00",x"00"),
  1599 => (x"00",x"00",x"00",x"00"),
  1600 => (x"00",x"12",x"64",x"00"),
  1601 => (x"00",x"2b",x"d2",x"00"),
  1602 => (x"00",x"00",x"00",x"00"),
  1603 => (x"00",x"00",x"12",x"64"),
  1604 => (x"00",x"00",x"2b",x"f0"),
  1605 => (x"64",x"00",x"00",x"00"),
  1606 => (x"00",x"00",x"00",x"12"),
  1607 => (x"00",x"00",x"00",x"00"),
  1608 => (x"12",x"f9",x"00",x"00"),
  1609 => (x"00",x"00",x"00",x"00"),
  1610 => (x"00",x"00",x"00",x"00"),
  1611 => (x"00",x"19",x"31",x"00"),
  1612 => (x"34",x"36",x"43",x"00"),
  1613 => (x"20",x"20",x"20",x"20"),
  1614 => (x"4d",x"4f",x"52",x"20"),
  1615 => (x"61",x"6f",x"4c",x"00"),
  1616 => (x"2e",x"2a",x"20",x"64"),
  1617 => (x"f0",x"fe",x"1e",x"00"),
  1618 => (x"cd",x"78",x"c0",x"48"),
  1619 => (x"26",x"09",x"79",x"09"),
  1620 => (x"fe",x"1e",x"1e",x"4f"),
  1621 => (x"48",x"7e",x"bf",x"f0"),
  1622 => (x"1e",x"4f",x"26",x"26"),
  1623 => (x"c1",x"48",x"f0",x"fe"),
  1624 => (x"1e",x"4f",x"26",x"78"),
  1625 => (x"c0",x"48",x"f0",x"fe"),
  1626 => (x"1e",x"4f",x"26",x"78"),
  1627 => (x"52",x"c0",x"4a",x"71"),
  1628 => (x"0e",x"4f",x"26",x"52"),
  1629 => (x"5d",x"5c",x"5b",x"5e"),
  1630 => (x"71",x"86",x"f4",x"0e"),
  1631 => (x"7e",x"6d",x"97",x"4d"),
  1632 => (x"97",x"4c",x"a5",x"c1"),
  1633 => (x"a6",x"c8",x"48",x"6c"),
  1634 => (x"c4",x"48",x"6e",x"58"),
  1635 => (x"c5",x"05",x"a8",x"66"),
  1636 => (x"c0",x"48",x"ff",x"87"),
  1637 => (x"ca",x"ff",x"87",x"e6"),
  1638 => (x"49",x"a5",x"c2",x"87"),
  1639 => (x"71",x"4b",x"6c",x"97"),
  1640 => (x"6b",x"97",x"4b",x"a3"),
  1641 => (x"7e",x"6c",x"97",x"4b"),
  1642 => (x"80",x"c1",x"48",x"6e"),
  1643 => (x"c7",x"58",x"a6",x"c8"),
  1644 => (x"58",x"a6",x"cc",x"98"),
  1645 => (x"fe",x"7c",x"97",x"70"),
  1646 => (x"48",x"73",x"87",x"e1"),
  1647 => (x"4d",x"26",x"8e",x"f4"),
  1648 => (x"4b",x"26",x"4c",x"26"),
  1649 => (x"5e",x"0e",x"4f",x"26"),
  1650 => (x"f4",x"0e",x"5c",x"5b"),
  1651 => (x"d8",x"4c",x"71",x"86"),
  1652 => (x"ff",x"c3",x"4a",x"66"),
  1653 => (x"4b",x"a4",x"c2",x"9a"),
  1654 => (x"73",x"49",x"6c",x"97"),
  1655 => (x"51",x"72",x"49",x"a1"),
  1656 => (x"6e",x"7e",x"6c",x"97"),
  1657 => (x"c8",x"80",x"c1",x"48"),
  1658 => (x"98",x"c7",x"58",x"a6"),
  1659 => (x"70",x"58",x"a6",x"cc"),
  1660 => (x"ff",x"8e",x"f4",x"54"),
  1661 => (x"1e",x"1e",x"87",x"ca"),
  1662 => (x"e0",x"87",x"e8",x"fd"),
  1663 => (x"c0",x"49",x"4a",x"bf"),
  1664 => (x"02",x"99",x"c0",x"e0"),
  1665 => (x"1e",x"72",x"87",x"cb"),
  1666 => (x"49",x"ce",x"f0",x"c2"),
  1667 => (x"c4",x"87",x"f7",x"fe"),
  1668 => (x"87",x"fd",x"fc",x"86"),
  1669 => (x"c2",x"fd",x"7e",x"70"),
  1670 => (x"4f",x"26",x"26",x"87"),
  1671 => (x"ce",x"f0",x"c2",x"1e"),
  1672 => (x"87",x"c7",x"fd",x"49"),
  1673 => (x"49",x"f6",x"e7",x"c1"),
  1674 => (x"c4",x"87",x"da",x"fc"),
  1675 => (x"4f",x"26",x"87",x"c8"),
  1676 => (x"48",x"d0",x"ff",x"1e"),
  1677 => (x"ff",x"78",x"e1",x"c8"),
  1678 => (x"78",x"c5",x"48",x"d4"),
  1679 => (x"c3",x"02",x"66",x"c4"),
  1680 => (x"78",x"e0",x"c3",x"87"),
  1681 => (x"c6",x"02",x"66",x"c8"),
  1682 => (x"48",x"d4",x"ff",x"87"),
  1683 => (x"ff",x"78",x"f0",x"c3"),
  1684 => (x"78",x"71",x"48",x"d4"),
  1685 => (x"c8",x"48",x"d0",x"ff"),
  1686 => (x"e0",x"c0",x"78",x"e1"),
  1687 => (x"0e",x"4f",x"26",x"78"),
  1688 => (x"0e",x"5c",x"5b",x"5e"),
  1689 => (x"f0",x"c2",x"4c",x"71"),
  1690 => (x"c6",x"fc",x"49",x"ce"),
  1691 => (x"c0",x"4a",x"70",x"87"),
  1692 => (x"c2",x"04",x"aa",x"b7"),
  1693 => (x"e0",x"c3",x"87",x"e3"),
  1694 => (x"87",x"c9",x"05",x"aa"),
  1695 => (x"48",x"e9",x"ec",x"c1"),
  1696 => (x"d4",x"c2",x"78",x"c1"),
  1697 => (x"aa",x"f0",x"c3",x"87"),
  1698 => (x"c1",x"87",x"c9",x"05"),
  1699 => (x"c1",x"48",x"e5",x"ec"),
  1700 => (x"87",x"f5",x"c1",x"78"),
  1701 => (x"bf",x"e9",x"ec",x"c1"),
  1702 => (x"72",x"87",x"c7",x"02"),
  1703 => (x"b3",x"c0",x"c2",x"4b"),
  1704 => (x"4b",x"72",x"87",x"c2"),
  1705 => (x"d1",x"05",x"9c",x"74"),
  1706 => (x"e5",x"ec",x"c1",x"87"),
  1707 => (x"ec",x"c1",x"1e",x"bf"),
  1708 => (x"72",x"1e",x"bf",x"e9"),
  1709 => (x"87",x"f8",x"fd",x"49"),
  1710 => (x"ec",x"c1",x"86",x"c8"),
  1711 => (x"c0",x"02",x"bf",x"e5"),
  1712 => (x"49",x"73",x"87",x"e0"),
  1713 => (x"91",x"29",x"b7",x"c4"),
  1714 => (x"81",x"c5",x"ee",x"c1"),
  1715 => (x"9a",x"cf",x"4a",x"73"),
  1716 => (x"48",x"c1",x"92",x"c2"),
  1717 => (x"4a",x"70",x"30",x"72"),
  1718 => (x"48",x"72",x"ba",x"ff"),
  1719 => (x"79",x"70",x"98",x"69"),
  1720 => (x"49",x"73",x"87",x"db"),
  1721 => (x"91",x"29",x"b7",x"c4"),
  1722 => (x"81",x"c5",x"ee",x"c1"),
  1723 => (x"9a",x"cf",x"4a",x"73"),
  1724 => (x"48",x"c3",x"92",x"c2"),
  1725 => (x"4a",x"70",x"30",x"72"),
  1726 => (x"70",x"b0",x"69",x"48"),
  1727 => (x"e9",x"ec",x"c1",x"79"),
  1728 => (x"c1",x"78",x"c0",x"48"),
  1729 => (x"c0",x"48",x"e5",x"ec"),
  1730 => (x"ce",x"f0",x"c2",x"78"),
  1731 => (x"87",x"e3",x"f9",x"49"),
  1732 => (x"b7",x"c0",x"4a",x"70"),
  1733 => (x"dd",x"fd",x"03",x"aa"),
  1734 => (x"c2",x"48",x"c0",x"87"),
  1735 => (x"26",x"4d",x"26",x"87"),
  1736 => (x"26",x"4b",x"26",x"4c"),
  1737 => (x"00",x"00",x"00",x"4f"),
  1738 => (x"00",x"00",x"00",x"00"),
  1739 => (x"4a",x"71",x"1e",x"00"),
  1740 => (x"87",x"eb",x"fc",x"49"),
  1741 => (x"c0",x"1e",x"4f",x"26"),
  1742 => (x"c4",x"49",x"72",x"4a"),
  1743 => (x"c5",x"ee",x"c1",x"91"),
  1744 => (x"c1",x"79",x"c0",x"81"),
  1745 => (x"aa",x"b7",x"d0",x"82"),
  1746 => (x"26",x"87",x"ee",x"04"),
  1747 => (x"5b",x"5e",x"0e",x"4f"),
  1748 => (x"71",x"0e",x"5d",x"5c"),
  1749 => (x"87",x"cb",x"f8",x"4d"),
  1750 => (x"b7",x"c4",x"4a",x"75"),
  1751 => (x"ee",x"c1",x"92",x"2a"),
  1752 => (x"4c",x"75",x"82",x"c5"),
  1753 => (x"94",x"c2",x"9c",x"cf"),
  1754 => (x"74",x"4b",x"49",x"6a"),
  1755 => (x"c2",x"9b",x"c3",x"2b"),
  1756 => (x"70",x"30",x"74",x"48"),
  1757 => (x"74",x"bc",x"ff",x"4c"),
  1758 => (x"70",x"98",x"71",x"48"),
  1759 => (x"87",x"db",x"f7",x"7a"),
  1760 => (x"d8",x"fe",x"48",x"73"),
  1761 => (x"00",x"00",x"00",x"87"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"00",x"00",x"00"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"00",x"00",x"00",x"00"),
  1776 => (x"00",x"00",x"00",x"00"),
  1777 => (x"d0",x"ff",x"1e",x"00"),
  1778 => (x"78",x"e1",x"c8",x"48"),
  1779 => (x"d4",x"ff",x"48",x"71"),
  1780 => (x"4f",x"26",x"78",x"08"),
  1781 => (x"48",x"d0",x"ff",x"1e"),
  1782 => (x"71",x"78",x"e1",x"c8"),
  1783 => (x"08",x"d4",x"ff",x"48"),
  1784 => (x"48",x"66",x"c4",x"78"),
  1785 => (x"78",x"08",x"d4",x"ff"),
  1786 => (x"71",x"1e",x"4f",x"26"),
  1787 => (x"49",x"66",x"c4",x"4a"),
  1788 => (x"ff",x"49",x"72",x"1e"),
  1789 => (x"d0",x"ff",x"87",x"de"),
  1790 => (x"78",x"e0",x"c0",x"48"),
  1791 => (x"1e",x"4f",x"26",x"26"),
  1792 => (x"4b",x"71",x"1e",x"73"),
  1793 => (x"1e",x"49",x"66",x"c8"),
  1794 => (x"e0",x"c1",x"4a",x"73"),
  1795 => (x"d9",x"ff",x"49",x"a2"),
  1796 => (x"87",x"c4",x"26",x"87"),
  1797 => (x"4c",x"26",x"4d",x"26"),
  1798 => (x"4f",x"26",x"4b",x"26"),
  1799 => (x"4a",x"d4",x"ff",x"1e"),
  1800 => (x"ff",x"7a",x"ff",x"c3"),
  1801 => (x"e1",x"c0",x"48",x"d0"),
  1802 => (x"c2",x"7a",x"de",x"78"),
  1803 => (x"7a",x"bf",x"d8",x"f0"),
  1804 => (x"28",x"c8",x"48",x"49"),
  1805 => (x"48",x"71",x"7a",x"70"),
  1806 => (x"7a",x"70",x"28",x"d0"),
  1807 => (x"28",x"d8",x"48",x"71"),
  1808 => (x"f0",x"c2",x"7a",x"70"),
  1809 => (x"49",x"7a",x"bf",x"dc"),
  1810 => (x"70",x"28",x"c8",x"48"),
  1811 => (x"d0",x"48",x"71",x"7a"),
  1812 => (x"71",x"7a",x"70",x"28"),
  1813 => (x"70",x"28",x"d8",x"48"),
  1814 => (x"48",x"d0",x"ff",x"7a"),
  1815 => (x"26",x"78",x"e0",x"c0"),
  1816 => (x"1e",x"73",x"1e",x"4f"),
  1817 => (x"f0",x"c2",x"4a",x"71"),
  1818 => (x"72",x"4b",x"bf",x"d8"),
  1819 => (x"aa",x"e0",x"c0",x"2b"),
  1820 => (x"72",x"87",x"ce",x"04"),
  1821 => (x"89",x"e0",x"c0",x"49"),
  1822 => (x"bf",x"dc",x"f0",x"c2"),
  1823 => (x"cf",x"2b",x"71",x"4b"),
  1824 => (x"49",x"e0",x"c0",x"87"),
  1825 => (x"f0",x"c2",x"89",x"72"),
  1826 => (x"71",x"48",x"bf",x"dc"),
  1827 => (x"b3",x"49",x"70",x"30"),
  1828 => (x"73",x"9b",x"66",x"c8"),
  1829 => (x"26",x"87",x"c4",x"48"),
  1830 => (x"26",x"4c",x"26",x"4d"),
  1831 => (x"0e",x"4f",x"26",x"4b"),
  1832 => (x"5d",x"5c",x"5b",x"5e"),
  1833 => (x"71",x"86",x"ec",x"0e"),
  1834 => (x"d8",x"f0",x"c2",x"4b"),
  1835 => (x"73",x"4c",x"7e",x"bf"),
  1836 => (x"ab",x"e0",x"c0",x"2c"),
  1837 => (x"87",x"e0",x"c0",x"04"),
  1838 => (x"c0",x"48",x"a6",x"c4"),
  1839 => (x"c0",x"49",x"73",x"78"),
  1840 => (x"4a",x"71",x"89",x"e0"),
  1841 => (x"48",x"66",x"e4",x"c0"),
  1842 => (x"a6",x"cc",x"30",x"72"),
  1843 => (x"dc",x"f0",x"c2",x"58"),
  1844 => (x"71",x"4c",x"4d",x"bf"),
  1845 => (x"87",x"e4",x"c0",x"2c"),
  1846 => (x"e4",x"c0",x"49",x"73"),
  1847 => (x"30",x"71",x"48",x"66"),
  1848 => (x"c0",x"58",x"a6",x"c8"),
  1849 => (x"89",x"73",x"49",x"e0"),
  1850 => (x"48",x"66",x"e4",x"c0"),
  1851 => (x"a6",x"cc",x"28",x"71"),
  1852 => (x"dc",x"f0",x"c2",x"58"),
  1853 => (x"71",x"48",x"4d",x"bf"),
  1854 => (x"b4",x"49",x"70",x"30"),
  1855 => (x"9c",x"66",x"e4",x"c0"),
  1856 => (x"e8",x"c0",x"84",x"c1"),
  1857 => (x"c2",x"04",x"ac",x"66"),
  1858 => (x"c0",x"4c",x"c0",x"87"),
  1859 => (x"d3",x"04",x"ab",x"e0"),
  1860 => (x"48",x"a6",x"cc",x"87"),
  1861 => (x"49",x"73",x"78",x"c0"),
  1862 => (x"74",x"89",x"e0",x"c0"),
  1863 => (x"d4",x"30",x"71",x"48"),
  1864 => (x"87",x"d5",x"58",x"a6"),
  1865 => (x"48",x"74",x"49",x"73"),
  1866 => (x"a6",x"d0",x"30",x"71"),
  1867 => (x"49",x"e0",x"c0",x"58"),
  1868 => (x"48",x"74",x"89",x"73"),
  1869 => (x"a6",x"d4",x"28",x"71"),
  1870 => (x"4a",x"66",x"c4",x"58"),
  1871 => (x"9a",x"6e",x"ba",x"ff"),
  1872 => (x"ff",x"49",x"66",x"c8"),
  1873 => (x"72",x"99",x"75",x"b9"),
  1874 => (x"b0",x"66",x"cc",x"48"),
  1875 => (x"58",x"dc",x"f0",x"c2"),
  1876 => (x"66",x"d0",x"48",x"71"),
  1877 => (x"e0",x"f0",x"c2",x"b0"),
  1878 => (x"87",x"c0",x"fb",x"58"),
  1879 => (x"f6",x"fc",x"8e",x"ec"),
  1880 => (x"d0",x"ff",x"1e",x"87"),
  1881 => (x"78",x"c9",x"c8",x"48"),
  1882 => (x"d4",x"ff",x"48",x"71"),
  1883 => (x"4f",x"26",x"78",x"08"),
  1884 => (x"49",x"4a",x"71",x"1e"),
  1885 => (x"d0",x"ff",x"87",x"eb"),
  1886 => (x"26",x"78",x"c8",x"48"),
  1887 => (x"1e",x"73",x"1e",x"4f"),
  1888 => (x"f0",x"c2",x"4b",x"71"),
  1889 => (x"c3",x"02",x"bf",x"ec"),
  1890 => (x"87",x"eb",x"c2",x"87"),
  1891 => (x"c8",x"48",x"d0",x"ff"),
  1892 => (x"49",x"73",x"78",x"c9"),
  1893 => (x"ff",x"b1",x"e0",x"c0"),
  1894 => (x"78",x"71",x"48",x"d4"),
  1895 => (x"48",x"e0",x"f0",x"c2"),
  1896 => (x"66",x"c8",x"78",x"c0"),
  1897 => (x"c3",x"87",x"c5",x"02"),
  1898 => (x"87",x"c2",x"49",x"ff"),
  1899 => (x"f0",x"c2",x"49",x"c0"),
  1900 => (x"66",x"cc",x"59",x"e8"),
  1901 => (x"c5",x"87",x"c6",x"02"),
  1902 => (x"c4",x"4a",x"d5",x"d5"),
  1903 => (x"ff",x"ff",x"cf",x"87"),
  1904 => (x"ec",x"f0",x"c2",x"4a"),
  1905 => (x"ec",x"f0",x"c2",x"5a"),
  1906 => (x"c4",x"78",x"c1",x"48"),
  1907 => (x"26",x"4d",x"26",x"87"),
  1908 => (x"26",x"4b",x"26",x"4c"),
  1909 => (x"5b",x"5e",x"0e",x"4f"),
  1910 => (x"71",x"0e",x"5d",x"5c"),
  1911 => (x"e8",x"f0",x"c2",x"4a"),
  1912 => (x"9a",x"72",x"4c",x"bf"),
  1913 => (x"49",x"87",x"cb",x"02"),
  1914 => (x"f5",x"c1",x"91",x"c8"),
  1915 => (x"83",x"71",x"4b",x"f3"),
  1916 => (x"f9",x"c1",x"87",x"c4"),
  1917 => (x"4d",x"c0",x"4b",x"f3"),
  1918 => (x"99",x"74",x"49",x"13"),
  1919 => (x"bf",x"e4",x"f0",x"c2"),
  1920 => (x"48",x"d4",x"ff",x"b9"),
  1921 => (x"b7",x"c1",x"78",x"71"),
  1922 => (x"b7",x"c8",x"85",x"2c"),
  1923 => (x"87",x"e8",x"04",x"ad"),
  1924 => (x"bf",x"e0",x"f0",x"c2"),
  1925 => (x"c2",x"80",x"c8",x"48"),
  1926 => (x"fe",x"58",x"e4",x"f0"),
  1927 => (x"73",x"1e",x"87",x"ef"),
  1928 => (x"13",x"4b",x"71",x"1e"),
  1929 => (x"cb",x"02",x"9a",x"4a"),
  1930 => (x"fe",x"49",x"72",x"87"),
  1931 => (x"4a",x"13",x"87",x"e7"),
  1932 => (x"87",x"f5",x"05",x"9a"),
  1933 => (x"1e",x"87",x"da",x"fe"),
  1934 => (x"bf",x"e0",x"f0",x"c2"),
  1935 => (x"e0",x"f0",x"c2",x"49"),
  1936 => (x"78",x"a1",x"c1",x"48"),
  1937 => (x"a9",x"b7",x"c0",x"c4"),
  1938 => (x"ff",x"87",x"db",x"03"),
  1939 => (x"f0",x"c2",x"48",x"d4"),
  1940 => (x"c2",x"78",x"bf",x"e4"),
  1941 => (x"49",x"bf",x"e0",x"f0"),
  1942 => (x"48",x"e0",x"f0",x"c2"),
  1943 => (x"c4",x"78",x"a1",x"c1"),
  1944 => (x"04",x"a9",x"b7",x"c0"),
  1945 => (x"d0",x"ff",x"87",x"e5"),
  1946 => (x"c2",x"78",x"c8",x"48"),
  1947 => (x"c0",x"48",x"ec",x"f0"),
  1948 => (x"00",x"4f",x"26",x"78"),
  1949 => (x"00",x"00",x"00",x"00"),
  1950 => (x"00",x"00",x"00",x"00"),
  1951 => (x"5f",x"5f",x"00",x"00"),
  1952 => (x"00",x"00",x"00",x"00"),
  1953 => (x"03",x"00",x"03",x"03"),
  1954 => (x"14",x"00",x"00",x"03"),
  1955 => (x"7f",x"14",x"7f",x"7f"),
  1956 => (x"00",x"00",x"14",x"7f"),
  1957 => (x"6b",x"6b",x"2e",x"24"),
  1958 => (x"4c",x"00",x"12",x"3a"),
  1959 => (x"6c",x"18",x"36",x"6a"),
  1960 => (x"30",x"00",x"32",x"56"),
  1961 => (x"77",x"59",x"4f",x"7e"),
  1962 => (x"00",x"40",x"68",x"3a"),
  1963 => (x"03",x"07",x"04",x"00"),
  1964 => (x"00",x"00",x"00",x"00"),
  1965 => (x"63",x"3e",x"1c",x"00"),
  1966 => (x"00",x"00",x"00",x"41"),
  1967 => (x"3e",x"63",x"41",x"00"),
  1968 => (x"08",x"00",x"00",x"1c"),
  1969 => (x"1c",x"1c",x"3e",x"2a"),
  1970 => (x"00",x"08",x"2a",x"3e"),
  1971 => (x"3e",x"3e",x"08",x"08"),
  1972 => (x"00",x"00",x"08",x"08"),
  1973 => (x"60",x"e0",x"80",x"00"),
  1974 => (x"00",x"00",x"00",x"00"),
  1975 => (x"08",x"08",x"08",x"08"),
  1976 => (x"00",x"00",x"08",x"08"),
  1977 => (x"60",x"60",x"00",x"00"),
  1978 => (x"40",x"00",x"00",x"00"),
  1979 => (x"0c",x"18",x"30",x"60"),
  1980 => (x"00",x"01",x"03",x"06"),
  1981 => (x"4d",x"59",x"7f",x"3e"),
  1982 => (x"00",x"00",x"3e",x"7f"),
  1983 => (x"7f",x"7f",x"06",x"04"),
  1984 => (x"00",x"00",x"00",x"00"),
  1985 => (x"59",x"71",x"63",x"42"),
  1986 => (x"00",x"00",x"46",x"4f"),
  1987 => (x"49",x"49",x"63",x"22"),
  1988 => (x"18",x"00",x"36",x"7f"),
  1989 => (x"7f",x"13",x"16",x"1c"),
  1990 => (x"00",x"00",x"10",x"7f"),
  1991 => (x"45",x"45",x"67",x"27"),
  1992 => (x"00",x"00",x"39",x"7d"),
  1993 => (x"49",x"4b",x"7e",x"3c"),
  1994 => (x"00",x"00",x"30",x"79"),
  1995 => (x"79",x"71",x"01",x"01"),
  1996 => (x"00",x"00",x"07",x"0f"),
  1997 => (x"49",x"49",x"7f",x"36"),
  1998 => (x"00",x"00",x"36",x"7f"),
  1999 => (x"69",x"49",x"4f",x"06"),
  2000 => (x"00",x"00",x"1e",x"3f"),
  2001 => (x"66",x"66",x"00",x"00"),
  2002 => (x"00",x"00",x"00",x"00"),
  2003 => (x"66",x"e6",x"80",x"00"),
  2004 => (x"00",x"00",x"00",x"00"),
  2005 => (x"14",x"14",x"08",x"08"),
  2006 => (x"00",x"00",x"22",x"22"),
  2007 => (x"14",x"14",x"14",x"14"),
  2008 => (x"00",x"00",x"14",x"14"),
  2009 => (x"14",x"14",x"22",x"22"),
  2010 => (x"00",x"00",x"08",x"08"),
  2011 => (x"59",x"51",x"03",x"02"),
  2012 => (x"3e",x"00",x"06",x"0f"),
  2013 => (x"55",x"5d",x"41",x"7f"),
  2014 => (x"00",x"00",x"1e",x"1f"),
  2015 => (x"09",x"09",x"7f",x"7e"),
  2016 => (x"00",x"00",x"7e",x"7f"),
  2017 => (x"49",x"49",x"7f",x"7f"),
  2018 => (x"00",x"00",x"36",x"7f"),
  2019 => (x"41",x"63",x"3e",x"1c"),
  2020 => (x"00",x"00",x"41",x"41"),
  2021 => (x"63",x"41",x"7f",x"7f"),
  2022 => (x"00",x"00",x"1c",x"3e"),
  2023 => (x"49",x"49",x"7f",x"7f"),
  2024 => (x"00",x"00",x"41",x"41"),
  2025 => (x"09",x"09",x"7f",x"7f"),
  2026 => (x"00",x"00",x"01",x"01"),
  2027 => (x"49",x"41",x"7f",x"3e"),
  2028 => (x"00",x"00",x"7a",x"7b"),
  2029 => (x"08",x"08",x"7f",x"7f"),
  2030 => (x"00",x"00",x"7f",x"7f"),
  2031 => (x"7f",x"7f",x"41",x"00"),
  2032 => (x"00",x"00",x"00",x"41"),
  2033 => (x"40",x"40",x"60",x"20"),
  2034 => (x"7f",x"00",x"3f",x"7f"),
  2035 => (x"36",x"1c",x"08",x"7f"),
  2036 => (x"00",x"00",x"41",x"63"),
  2037 => (x"40",x"40",x"7f",x"7f"),
  2038 => (x"7f",x"00",x"40",x"40"),
  2039 => (x"06",x"0c",x"06",x"7f"),
  2040 => (x"7f",x"00",x"7f",x"7f"),
  2041 => (x"18",x"0c",x"06",x"7f"),
  2042 => (x"00",x"00",x"7f",x"7f"),
  2043 => (x"41",x"41",x"7f",x"3e"),
  2044 => (x"00",x"00",x"3e",x"7f"),
  2045 => (x"09",x"09",x"7f",x"7f"),
  2046 => (x"3e",x"00",x"06",x"0f"),
  2047 => (x"7f",x"61",x"41",x"7f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

