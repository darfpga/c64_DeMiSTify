library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f0f1c287",
    12 => x"86c0c64e",
    13 => x"49f0f1c2",
    14 => x"48f8dec2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087d9e1",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"4a711e4f",
    50 => x"484966c4",
    51 => x"a6c888c1",
    52 => x"02997158",
    53 => x"481287d4",
    54 => x"7808d4ff",
    55 => x"484966c4",
    56 => x"a6c888c1",
    57 => x"05997158",
    58 => x"4f2687ec",
    59 => x"c44a711e",
    60 => x"c1484966",
    61 => x"58a6c888",
    62 => x"d6029971",
    63 => x"48d4ff87",
    64 => x"6878ffc3",
    65 => x"4966c452",
    66 => x"c888c148",
    67 => x"997158a6",
    68 => x"2687ea05",
    69 => x"1e731e4f",
    70 => x"c34bd4ff",
    71 => x"4a6b7bff",
    72 => x"6b7bffc3",
    73 => x"7232c849",
    74 => x"7bffc3b1",
    75 => x"31c84a6b",
    76 => x"ffc3b271",
    77 => x"c8496b7b",
    78 => x"71b17232",
    79 => x"2687c448",
    80 => x"264c264d",
    81 => x"0e4f264b",
    82 => x"5d5c5b5e",
    83 => x"ff4a710e",
    84 => x"49724cd4",
    85 => x"7199ffc3",
    86 => x"f8dec27c",
    87 => x"87c805bf",
    88 => x"c94866d0",
    89 => x"58a6d430",
    90 => x"d84966d0",
    91 => x"99ffc329",
    92 => x"66d07c71",
    93 => x"c329d049",
    94 => x"7c7199ff",
    95 => x"c84966d0",
    96 => x"99ffc329",
    97 => x"66d07c71",
    98 => x"99ffc349",
    99 => x"49727c71",
   100 => x"ffc329d0",
   101 => x"6c7c7199",
   102 => x"fff0c94b",
   103 => x"abffc34d",
   104 => x"c387d005",
   105 => x"4b6c7cff",
   106 => x"c6028dc1",
   107 => x"abffc387",
   108 => x"7387f002",
   109 => x"87c7fe48",
   110 => x"ff49c01e",
   111 => x"ffc348d4",
   112 => x"c381c178",
   113 => x"04a9b7c8",
   114 => x"4f2687f1",
   115 => x"e71e731e",
   116 => x"dff8c487",
   117 => x"c01ec04b",
   118 => x"f7c1f0ff",
   119 => x"87e7fd49",
   120 => x"a8c186c4",
   121 => x"87eac005",
   122 => x"c348d4ff",
   123 => x"c0c178ff",
   124 => x"c0c0c0c0",
   125 => x"f0e1c01e",
   126 => x"fd49e9c1",
   127 => x"86c487c9",
   128 => x"ca059870",
   129 => x"48d4ff87",
   130 => x"c178ffc3",
   131 => x"fe87cb48",
   132 => x"8bc187e6",
   133 => x"87fdfe05",
   134 => x"e6fc48c0",
   135 => x"1e731e87",
   136 => x"c348d4ff",
   137 => x"4bd378ff",
   138 => x"ffc01ec0",
   139 => x"49c1c1f0",
   140 => x"c487d4fc",
   141 => x"05987086",
   142 => x"d4ff87ca",
   143 => x"78ffc348",
   144 => x"87cb48c1",
   145 => x"c187f1fd",
   146 => x"dbff058b",
   147 => x"fb48c087",
   148 => x"5e0e87f1",
   149 => x"ff0e5c5b",
   150 => x"dbfd4cd4",
   151 => x"1eeac687",
   152 => x"c1f0e1c0",
   153 => x"defb49c8",
   154 => x"c186c487",
   155 => x"87c802a8",
   156 => x"c087eafe",
   157 => x"87e2c148",
   158 => x"7087dafa",
   159 => x"ffffcf49",
   160 => x"a9eac699",
   161 => x"fe87c802",
   162 => x"48c087d3",
   163 => x"c387cbc1",
   164 => x"f1c07cff",
   165 => x"87f4fc4b",
   166 => x"c0029870",
   167 => x"1ec087eb",
   168 => x"c1f0ffc0",
   169 => x"defa49fa",
   170 => x"7086c487",
   171 => x"87d90598",
   172 => x"6c7cffc3",
   173 => x"7cffc349",
   174 => x"c17c7c7c",
   175 => x"c40299c0",
   176 => x"d548c187",
   177 => x"d148c087",
   178 => x"05abc287",
   179 => x"48c087c4",
   180 => x"8bc187c8",
   181 => x"87fdfe05",
   182 => x"e4f948c0",
   183 => x"1e731e87",
   184 => x"48f8dec2",
   185 => x"4bc778c1",
   186 => x"c248d0ff",
   187 => x"87c8fb78",
   188 => x"c348d0ff",
   189 => x"c01ec078",
   190 => x"c0c1d0e5",
   191 => x"87c7f949",
   192 => x"a8c186c4",
   193 => x"4b87c105",
   194 => x"c505abc2",
   195 => x"c048c087",
   196 => x"8bc187f9",
   197 => x"87d0ff05",
   198 => x"c287f7fc",
   199 => x"7058fcde",
   200 => x"87cd0598",
   201 => x"ffc01ec1",
   202 => x"49d0c1f0",
   203 => x"c487d8f8",
   204 => x"48d4ff86",
   205 => x"c478ffc3",
   206 => x"dfc287de",
   207 => x"d0ff58c0",
   208 => x"ff78c248",
   209 => x"ffc348d4",
   210 => x"f748c178",
   211 => x"5e0e87f5",
   212 => x"0e5d5c5b",
   213 => x"ffc34a71",
   214 => x"4cd4ff4d",
   215 => x"d0ff7c75",
   216 => x"78c3c448",
   217 => x"1e727c75",
   218 => x"c1f0ffc0",
   219 => x"d6f749d8",
   220 => x"7086c487",
   221 => x"87c50298",
   222 => x"f0c048c1",
   223 => x"c37c7587",
   224 => x"c0c87cfe",
   225 => x"4966d41e",
   226 => x"c487faf4",
   227 => x"757c7586",
   228 => x"d87c757c",
   229 => x"754be0da",
   230 => x"99496c7c",
   231 => x"c187c505",
   232 => x"87f3058b",
   233 => x"d0ff7c75",
   234 => x"c078c248",
   235 => x"87cff648",
   236 => x"5c5b5e0e",
   237 => x"4b710e5d",
   238 => x"eec54cc0",
   239 => x"ff4adfcd",
   240 => x"ffc348d4",
   241 => x"c3496878",
   242 => x"c005a9fe",
   243 => x"4d7087fd",
   244 => x"cc029b73",
   245 => x"1e66d087",
   246 => x"cff44973",
   247 => x"d686c487",
   248 => x"48d0ff87",
   249 => x"c378d1c4",
   250 => x"66d07dff",
   251 => x"d488c148",
   252 => x"987058a6",
   253 => x"ff87f005",
   254 => x"ffc348d4",
   255 => x"9b737878",
   256 => x"ff87c505",
   257 => x"78d048d0",
   258 => x"c14c4ac1",
   259 => x"eefe058a",
   260 => x"f4487487",
   261 => x"731e87e9",
   262 => x"c04a711e",
   263 => x"48d4ff4b",
   264 => x"ff78ffc3",
   265 => x"c3c448d0",
   266 => x"48d4ff78",
   267 => x"7278ffc3",
   268 => x"f0ffc01e",
   269 => x"f449d1c1",
   270 => x"86c487cd",
   271 => x"d2059870",
   272 => x"1ec0c887",
   273 => x"fd4966cc",
   274 => x"86c487e6",
   275 => x"d0ff4b70",
   276 => x"7378c248",
   277 => x"87ebf348",
   278 => x"5c5b5e0e",
   279 => x"1ec00e5d",
   280 => x"c1f0ffc0",
   281 => x"def349c9",
   282 => x"c21ed287",
   283 => x"fc49c0df",
   284 => x"86c887fe",
   285 => x"84c14cc0",
   286 => x"04acb7d2",
   287 => x"dfc287f8",
   288 => x"49bf97c0",
   289 => x"c199c0c3",
   290 => x"c005a9c0",
   291 => x"dfc287e7",
   292 => x"49bf97c7",
   293 => x"dfc231d0",
   294 => x"4abf97c8",
   295 => x"b17232c8",
   296 => x"97c9dfc2",
   297 => x"71b14abf",
   298 => x"ffffcf4c",
   299 => x"84c19cff",
   300 => x"e7c134ca",
   301 => x"c9dfc287",
   302 => x"c149bf97",
   303 => x"c299c631",
   304 => x"bf97cadf",
   305 => x"2ab7c74a",
   306 => x"dfc2b172",
   307 => x"4abf97c5",
   308 => x"c29dcf4d",
   309 => x"bf97c6df",
   310 => x"ca9ac34a",
   311 => x"c7dfc232",
   312 => x"c24bbf97",
   313 => x"c2b27333",
   314 => x"bf97c8df",
   315 => x"9bc0c34b",
   316 => x"732bb7c6",
   317 => x"c181c2b2",
   318 => x"70307148",
   319 => x"7548c149",
   320 => x"724d7030",
   321 => x"7184c14c",
   322 => x"b7c0c894",
   323 => x"87cc06ad",
   324 => x"2db734c1",
   325 => x"adb7c0c8",
   326 => x"87f4ff01",
   327 => x"def04874",
   328 => x"5b5e0e87",
   329 => x"f80e5d5c",
   330 => x"e6e7c286",
   331 => x"c278c048",
   332 => x"c01ededf",
   333 => x"87defb49",
   334 => x"987086c4",
   335 => x"c087c505",
   336 => x"87cec948",
   337 => x"7ec14dc0",
   338 => x"bfc0f3c0",
   339 => x"d4e0c249",
   340 => x"4bc8714a",
   341 => x"7087d3ec",
   342 => x"87c20598",
   343 => x"f2c07ec0",
   344 => x"c249bffc",
   345 => x"714af0e0",
   346 => x"fdeb4bc8",
   347 => x"05987087",
   348 => x"7ec087c2",
   349 => x"fdc0026e",
   350 => x"e4e6c287",
   351 => x"e7c24dbf",
   352 => x"7ebf9fdc",
   353 => x"ead6c548",
   354 => x"87c705a8",
   355 => x"bfe4e6c2",
   356 => x"6e87ce4d",
   357 => x"d5e9ca48",
   358 => x"87c502a8",
   359 => x"f1c748c0",
   360 => x"dedfc287",
   361 => x"f949751e",
   362 => x"86c487ec",
   363 => x"c5059870",
   364 => x"c748c087",
   365 => x"f2c087dc",
   366 => x"c249bffc",
   367 => x"714af0e0",
   368 => x"e5ea4bc8",
   369 => x"05987087",
   370 => x"e7c287c8",
   371 => x"78c148e6",
   372 => x"f3c087da",
   373 => x"c249bfc0",
   374 => x"714ad4e0",
   375 => x"c9ea4bc8",
   376 => x"02987087",
   377 => x"c087c5c0",
   378 => x"87e6c648",
   379 => x"97dce7c2",
   380 => x"d5c149bf",
   381 => x"cdc005a9",
   382 => x"dde7c287",
   383 => x"c249bf97",
   384 => x"c002a9ea",
   385 => x"48c087c5",
   386 => x"c287c7c6",
   387 => x"bf97dedf",
   388 => x"e9c3487e",
   389 => x"cec002a8",
   390 => x"c3486e87",
   391 => x"c002a8eb",
   392 => x"48c087c5",
   393 => x"c287ebc5",
   394 => x"bf97e9df",
   395 => x"c0059949",
   396 => x"dfc287cc",
   397 => x"49bf97ea",
   398 => x"c002a9c2",
   399 => x"48c087c5",
   400 => x"c287cfc5",
   401 => x"bf97ebdf",
   402 => x"e2e7c248",
   403 => x"484c7058",
   404 => x"e7c288c1",
   405 => x"dfc258e6",
   406 => x"49bf97ec",
   407 => x"dfc28175",
   408 => x"4abf97ed",
   409 => x"a17232c8",
   410 => x"f3ebc27e",
   411 => x"c2786e48",
   412 => x"bf97eedf",
   413 => x"58a6c848",
   414 => x"bfe6e7c2",
   415 => x"87d4c202",
   416 => x"bffcf2c0",
   417 => x"f0e0c249",
   418 => x"4bc8714a",
   419 => x"7087dbe7",
   420 => x"c5c00298",
   421 => x"c348c087",
   422 => x"e7c287f8",
   423 => x"c24cbfde",
   424 => x"c25cc7ec",
   425 => x"bf97c3e0",
   426 => x"c231c849",
   427 => x"bf97c2e0",
   428 => x"c249a14a",
   429 => x"bf97c4e0",
   430 => x"7232d04a",
   431 => x"e0c249a1",
   432 => x"4abf97c5",
   433 => x"a17232d8",
   434 => x"9166c449",
   435 => x"bff3ebc2",
   436 => x"fbebc281",
   437 => x"cbe0c259",
   438 => x"c84abf97",
   439 => x"cae0c232",
   440 => x"a24bbf97",
   441 => x"cce0c24a",
   442 => x"d04bbf97",
   443 => x"4aa27333",
   444 => x"97cde0c2",
   445 => x"9bcf4bbf",
   446 => x"a27333d8",
   447 => x"ffebc24a",
   448 => x"fbebc25a",
   449 => x"8ac24abf",
   450 => x"ebc29274",
   451 => x"a17248ff",
   452 => x"87cac178",
   453 => x"97f0dfc2",
   454 => x"31c849bf",
   455 => x"97efdfc2",
   456 => x"49a14abf",
   457 => x"59eee7c2",
   458 => x"bfeae7c2",
   459 => x"c731c549",
   460 => x"29c981ff",
   461 => x"59c7ecc2",
   462 => x"97f5dfc2",
   463 => x"32c84abf",
   464 => x"97f4dfc2",
   465 => x"4aa24bbf",
   466 => x"6e9266c4",
   467 => x"c3ecc282",
   468 => x"fbebc25a",
   469 => x"c278c048",
   470 => x"7248f7eb",
   471 => x"ecc278a1",
   472 => x"ebc248c7",
   473 => x"c278bffb",
   474 => x"c248cbec",
   475 => x"78bfffeb",
   476 => x"bfe6e7c2",
   477 => x"87c9c002",
   478 => x"30c44874",
   479 => x"c9c07e70",
   480 => x"c3ecc287",
   481 => x"30c448bf",
   482 => x"e7c27e70",
   483 => x"786e48ea",
   484 => x"8ef848c1",
   485 => x"4c264d26",
   486 => x"4f264b26",
   487 => x"5c5b5e0e",
   488 => x"4a710e5d",
   489 => x"bfe6e7c2",
   490 => x"7287cb02",
   491 => x"722bc74b",
   492 => x"9cffc14c",
   493 => x"4b7287c9",
   494 => x"4c722bc8",
   495 => x"c29cffc3",
   496 => x"83bff3eb",
   497 => x"bff8f2c0",
   498 => x"87d902ab",
   499 => x"5bfcf2c0",
   500 => x"1ededfc2",
   501 => x"fdf04973",
   502 => x"7086c487",
   503 => x"87c50598",
   504 => x"e6c048c0",
   505 => x"e6e7c287",
   506 => x"87d202bf",
   507 => x"91c44974",
   508 => x"81dedfc2",
   509 => x"ffcf4d69",
   510 => x"9dffffff",
   511 => x"497487cb",
   512 => x"dfc291c2",
   513 => x"699f81de",
   514 => x"fe48754d",
   515 => x"5e0e87c6",
   516 => x"0e5d5c5b",
   517 => x"4c7186f8",
   518 => x"87c5059c",
   519 => x"c2c348c0",
   520 => x"7ea4c887",
   521 => x"78c0486e",
   522 => x"c70266d8",
   523 => x"9766d887",
   524 => x"87c505bf",
   525 => x"eac248c0",
   526 => x"c11ec087",
   527 => x"87ddca49",
   528 => x"4d7086c4",
   529 => x"c3c1029d",
   530 => x"eee7c287",
   531 => x"4966d84a",
   532 => x"87fbdfff",
   533 => x"c0029870",
   534 => x"4a7587f2",
   535 => x"cb4966d8",
   536 => x"87e0e04b",
   537 => x"c0029870",
   538 => x"1ec087e2",
   539 => x"c7029d75",
   540 => x"48a6c887",
   541 => x"87c578c0",
   542 => x"c148a6c8",
   543 => x"4966c878",
   544 => x"c487dac9",
   545 => x"9d4d7086",
   546 => x"87fdfe05",
   547 => x"c1029d75",
   548 => x"a5dc87cf",
   549 => x"69486e49",
   550 => x"49a5da78",
   551 => x"c448a6c4",
   552 => x"699f78a4",
   553 => x"0866c448",
   554 => x"e6e7c278",
   555 => x"87d202bf",
   556 => x"9f49a5d4",
   557 => x"ffc04969",
   558 => x"487199ff",
   559 => x"7e7030d0",
   560 => x"7ec087c2",
   561 => x"c448496e",
   562 => x"c480bf66",
   563 => x"c0780866",
   564 => x"49a4cc7c",
   565 => x"79bf66c4",
   566 => x"c049a4d0",
   567 => x"c248c179",
   568 => x"f848c087",
   569 => x"87ecfa8e",
   570 => x"5c5b5e0e",
   571 => x"4c710e5d",
   572 => x"cac1029c",
   573 => x"49a4c887",
   574 => x"c2c10269",
   575 => x"4a66d087",
   576 => x"d482496c",
   577 => x"66d05aa6",
   578 => x"e7c2b94d",
   579 => x"ff4abfe2",
   580 => x"719972ba",
   581 => x"e4c00299",
   582 => x"4ba4c487",
   583 => x"fbf9496b",
   584 => x"c27b7087",
   585 => x"49bfdee7",
   586 => x"7c71816c",
   587 => x"e7c2b975",
   588 => x"ff4abfe2",
   589 => x"719972ba",
   590 => x"dcff0599",
   591 => x"f97c7587",
   592 => x"731e87d2",
   593 => x"9b4b711e",
   594 => x"c887c702",
   595 => x"056949a3",
   596 => x"48c087c5",
   597 => x"c287f7c0",
   598 => x"4abff7eb",
   599 => x"6949a3c4",
   600 => x"c289c249",
   601 => x"91bfdee7",
   602 => x"c24aa271",
   603 => x"49bfe2e7",
   604 => x"a271996b",
   605 => x"fcf2c04a",
   606 => x"1e66c85a",
   607 => x"d5ea4972",
   608 => x"7086c487",
   609 => x"87c40598",
   610 => x"87c248c0",
   611 => x"c7f848c1",
   612 => x"1e731e87",
   613 => x"029b4b71",
   614 => x"a3c887c7",
   615 => x"c5056949",
   616 => x"c048c087",
   617 => x"ebc287f7",
   618 => x"c44abff7",
   619 => x"496949a3",
   620 => x"e7c289c2",
   621 => x"7191bfde",
   622 => x"e7c24aa2",
   623 => x"6b49bfe2",
   624 => x"4aa27199",
   625 => x"5afcf2c0",
   626 => x"721e66c8",
   627 => x"87fee549",
   628 => x"987086c4",
   629 => x"c087c405",
   630 => x"c187c248",
   631 => x"87f8f648",
   632 => x"5c5b5e0e",
   633 => x"711e0e5d",
   634 => x"4c66d44b",
   635 => x"9b732cc9",
   636 => x"87cfc102",
   637 => x"6949a3c8",
   638 => x"87c7c102",
   639 => x"d44da3d0",
   640 => x"e7c27d66",
   641 => x"ff49bfe2",
   642 => x"994a6bb9",
   643 => x"03ac717e",
   644 => x"7bc087cd",
   645 => x"4aa3cc7d",
   646 => x"6a49a3c4",
   647 => x"7287c279",
   648 => x"029c748c",
   649 => x"1e4987dd",
   650 => x"fbfa4973",
   651 => x"d486c487",
   652 => x"ffc74966",
   653 => x"87cb0299",
   654 => x"1ededfc2",
   655 => x"c1fc4973",
   656 => x"2686c487",
   657 => x"1e87cdf5",
   658 => x"4b711e73",
   659 => x"e4c0029b",
   660 => x"cbecc287",
   661 => x"c24a735b",
   662 => x"dee7c28a",
   663 => x"c29249bf",
   664 => x"48bff7eb",
   665 => x"ecc28072",
   666 => x"487158cf",
   667 => x"e7c230c4",
   668 => x"edc058ee",
   669 => x"c7ecc287",
   670 => x"fbebc248",
   671 => x"ecc278bf",
   672 => x"ebc248cb",
   673 => x"c278bfff",
   674 => x"02bfe6e7",
   675 => x"e7c287c9",
   676 => x"c449bfde",
   677 => x"c287c731",
   678 => x"49bfc3ec",
   679 => x"e7c231c4",
   680 => x"f3f359ee",
   681 => x"5b5e0e87",
   682 => x"4a710e5c",
   683 => x"9a724bc0",
   684 => x"87e1c002",
   685 => x"9f49a2da",
   686 => x"e7c24b69",
   687 => x"cf02bfe6",
   688 => x"49a2d487",
   689 => x"4c49699f",
   690 => x"9cffffc0",
   691 => x"87c234d0",
   692 => x"49744cc0",
   693 => x"fd4973b3",
   694 => x"f9f287ed",
   695 => x"5b5e0e87",
   696 => x"f40e5d5c",
   697 => x"c04a7186",
   698 => x"029a727e",
   699 => x"dfc287d8",
   700 => x"78c048da",
   701 => x"48d2dfc2",
   702 => x"bfcbecc2",
   703 => x"d6dfc278",
   704 => x"c7ecc248",
   705 => x"e7c278bf",
   706 => x"50c048fb",
   707 => x"bfeae7c2",
   708 => x"dadfc249",
   709 => x"aa714abf",
   710 => x"87c9c403",
   711 => x"99cf4972",
   712 => x"87e9c005",
   713 => x"48f8f2c0",
   714 => x"bfd2dfc2",
   715 => x"dedfc278",
   716 => x"d2dfc21e",
   717 => x"dfc249bf",
   718 => x"a1c148d2",
   719 => x"d5e37178",
   720 => x"c086c487",
   721 => x"c248f4f2",
   722 => x"cc78dedf",
   723 => x"f4f2c087",
   724 => x"e0c048bf",
   725 => x"f8f2c080",
   726 => x"dadfc258",
   727 => x"80c148bf",
   728 => x"58dedfc2",
   729 => x"000cb427",
   730 => x"bf97bf00",
   731 => x"c2029d4d",
   732 => x"e5c387e3",
   733 => x"dcc202ad",
   734 => x"f4f2c087",
   735 => x"a3cb4bbf",
   736 => x"cf4c1149",
   737 => x"d2c105ac",
   738 => x"df497587",
   739 => x"cd89c199",
   740 => x"eee7c291",
   741 => x"4aa3c181",
   742 => x"a3c35112",
   743 => x"c551124a",
   744 => x"51124aa3",
   745 => x"124aa3c7",
   746 => x"4aa3c951",
   747 => x"a3ce5112",
   748 => x"d051124a",
   749 => x"51124aa3",
   750 => x"124aa3d2",
   751 => x"4aa3d451",
   752 => x"a3d65112",
   753 => x"d851124a",
   754 => x"51124aa3",
   755 => x"124aa3dc",
   756 => x"4aa3de51",
   757 => x"7ec15112",
   758 => x"7487fac0",
   759 => x"0599c849",
   760 => x"7487ebc0",
   761 => x"0599d049",
   762 => x"66dc87d1",
   763 => x"87cbc002",
   764 => x"66dc4973",
   765 => x"0298700f",
   766 => x"6e87d3c0",
   767 => x"87c6c005",
   768 => x"48eee7c2",
   769 => x"f2c050c0",
   770 => x"c248bff4",
   771 => x"e7c287e1",
   772 => x"50c048fb",
   773 => x"eae7c27e",
   774 => x"dfc249bf",
   775 => x"714abfda",
   776 => x"f7fb04aa",
   777 => x"cbecc287",
   778 => x"c8c005bf",
   779 => x"e6e7c287",
   780 => x"f8c102bf",
   781 => x"d6dfc287",
   782 => x"dfed49bf",
   783 => x"c2497087",
   784 => x"c459dadf",
   785 => x"dfc248a6",
   786 => x"c278bfd6",
   787 => x"02bfe6e7",
   788 => x"c487d8c0",
   789 => x"ffcf4966",
   790 => x"99f8ffff",
   791 => x"c5c002a9",
   792 => x"c04cc087",
   793 => x"4cc187e1",
   794 => x"c487dcc0",
   795 => x"ffcf4966",
   796 => x"02a999f8",
   797 => x"c887c8c0",
   798 => x"78c048a6",
   799 => x"c887c5c0",
   800 => x"78c148a6",
   801 => x"744c66c8",
   802 => x"e0c0059c",
   803 => x"4966c487",
   804 => x"e7c289c2",
   805 => x"914abfde",
   806 => x"bff7ebc2",
   807 => x"d2dfc24a",
   808 => x"78a17248",
   809 => x"48dadfc2",
   810 => x"dff978c0",
   811 => x"f448c087",
   812 => x"87e0eb8e",
   813 => x"00000000",
   814 => x"ffffffff",
   815 => x"00000cc4",
   816 => x"00000ccd",
   817 => x"33544146",
   818 => x"20202032",
   819 => x"54414600",
   820 => x"20203631",
   821 => x"ff1e0020",
   822 => x"ffc348d4",
   823 => x"26486878",
   824 => x"d4ff1e4f",
   825 => x"78ffc348",
   826 => x"c048d0ff",
   827 => x"d4ff78e1",
   828 => x"c278d448",
   829 => x"ff48cfec",
   830 => x"2650bfd4",
   831 => x"d0ff1e4f",
   832 => x"78e0c048",
   833 => x"ff1e4f26",
   834 => x"497087cc",
   835 => x"87c60299",
   836 => x"05a9fbc0",
   837 => x"487187f1",
   838 => x"5e0e4f26",
   839 => x"710e5c5b",
   840 => x"fe4cc04b",
   841 => x"497087f0",
   842 => x"f9c00299",
   843 => x"a9ecc087",
   844 => x"87f2c002",
   845 => x"02a9fbc0",
   846 => x"cc87ebc0",
   847 => x"03acb766",
   848 => x"66d087c7",
   849 => x"7187c202",
   850 => x"02997153",
   851 => x"84c187c2",
   852 => x"7087c3fe",
   853 => x"cd029949",
   854 => x"a9ecc087",
   855 => x"c087c702",
   856 => x"ff05a9fb",
   857 => x"66d087d5",
   858 => x"c087c302",
   859 => x"ecc07b97",
   860 => x"87c405a9",
   861 => x"87c54a74",
   862 => x"0ac04a74",
   863 => x"c248728a",
   864 => x"264d2687",
   865 => x"264b264c",
   866 => x"c9fd1e4f",
   867 => x"c0497087",
   868 => x"04a9b7f0",
   869 => x"f9c087ca",
   870 => x"c301a9b7",
   871 => x"89f0c087",
   872 => x"a9b7c1c1",
   873 => x"c187ca04",
   874 => x"01a9b7da",
   875 => x"f7c087c3",
   876 => x"b7e1c189",
   877 => x"87ca04a9",
   878 => x"a9b7fac1",
   879 => x"c087c301",
   880 => x"487189fd",
   881 => x"5e0e4f26",
   882 => x"710e5c5b",
   883 => x"4cd4ff4a",
   884 => x"e9c04972",
   885 => x"9b4b7087",
   886 => x"c187c202",
   887 => x"48d0ff8b",
   888 => x"d5c178c5",
   889 => x"c649737c",
   890 => x"fae2c131",
   891 => x"484abf97",
   892 => x"7c70b071",
   893 => x"c448d0ff",
   894 => x"fe487378",
   895 => x"5e0e87c5",
   896 => x"0e5d5c5b",
   897 => x"4c7186f8",
   898 => x"d4fb7ec0",
   899 => x"c04bc087",
   900 => x"bf97ebfa",
   901 => x"04a9c049",
   902 => x"e9fb87cf",
   903 => x"c083c187",
   904 => x"bf97ebfa",
   905 => x"f106ab49",
   906 => x"ebfac087",
   907 => x"cf02bf97",
   908 => x"87e2fa87",
   909 => x"02994970",
   910 => x"ecc087c6",
   911 => x"87f105a9",
   912 => x"d1fa4bc0",
   913 => x"fa4d7087",
   914 => x"a6c887cc",
   915 => x"87c6fa58",
   916 => x"83c14a70",
   917 => x"9749a4c8",
   918 => x"02ad4969",
   919 => x"ffc087c7",
   920 => x"e7c005ad",
   921 => x"49a4c987",
   922 => x"c4496997",
   923 => x"c702a966",
   924 => x"ffc04887",
   925 => x"87d405a8",
   926 => x"9749a4ca",
   927 => x"02aa4969",
   928 => x"ffc087c6",
   929 => x"87c405aa",
   930 => x"87d07ec1",
   931 => x"02adecc0",
   932 => x"fbc087c6",
   933 => x"87c405ad",
   934 => x"7ec14bc0",
   935 => x"e1fe026e",
   936 => x"87d9f987",
   937 => x"8ef84873",
   938 => x"0087d6fb",
   939 => x"5c5b5e0e",
   940 => x"711e0e5d",
   941 => x"4bd4ff4d",
   942 => x"ecc21e75",
   943 => x"cde549d4",
   944 => x"7086c487",
   945 => x"d5c30298",
   946 => x"dcecc287",
   947 => x"49754cbf",
   948 => x"ff87f3fb",
   949 => x"78c548d0",
   950 => x"c07bd6c1",
   951 => x"49a2754a",
   952 => x"82c17b11",
   953 => x"04aab7cb",
   954 => x"4acc87f3",
   955 => x"c17bffc3",
   956 => x"b7e0c082",
   957 => x"87f404aa",
   958 => x"c448d0ff",
   959 => x"7bffc378",
   960 => x"d3c178c5",
   961 => x"c47bc17b",
   962 => x"029c7478",
   963 => x"c287ffc1",
   964 => x"c87ededf",
   965 => x"c08c4dc0",
   966 => x"c603acb7",
   967 => x"a4c0c887",
   968 => x"c84cc04d",
   969 => x"dc05adc0",
   970 => x"cfecc287",
   971 => x"d049bf97",
   972 => x"87d10299",
   973 => x"ecc21ec0",
   974 => x"c5e849d4",
   975 => x"7086c487",
   976 => x"eec04a49",
   977 => x"dedfc287",
   978 => x"d4ecc21e",
   979 => x"87f2e749",
   980 => x"497086c4",
   981 => x"48d0ff4a",
   982 => x"c178c5c8",
   983 => x"976e7bd4",
   984 => x"486e7bbf",
   985 => x"7e7080c1",
   986 => x"ff058dc1",
   987 => x"d0ff87f0",
   988 => x"7278c448",
   989 => x"87c5059a",
   990 => x"e3c048c0",
   991 => x"c21ec187",
   992 => x"e549d4ec",
   993 => x"86c487e2",
   994 => x"fe059c74",
   995 => x"d0ff87c1",
   996 => x"c178c548",
   997 => x"7bc07bd3",
   998 => x"48c178c4",
   999 => x"48c087c2",
  1000 => x"264d2626",
  1001 => x"264b264c",
  1002 => x"5b5e0e4f",
  1003 => x"1e0e5d5c",
  1004 => x"4cc04b71",
  1005 => x"c004ab4d",
  1006 => x"f7c087e8",
  1007 => x"9d751efe",
  1008 => x"c087c402",
  1009 => x"c187c24a",
  1010 => x"ec49724a",
  1011 => x"86c487cf",
  1012 => x"84c17e70",
  1013 => x"87c2056e",
  1014 => x"85c14c73",
  1015 => x"ff06ac73",
  1016 => x"486e87d8",
  1017 => x"87f9fe26",
  1018 => x"5c5b5e0e",
  1019 => x"cc4b710e",
  1020 => x"87d80266",
  1021 => x"8cf0c04c",
  1022 => x"7487d802",
  1023 => x"028ac14a",
  1024 => x"028a87d1",
  1025 => x"028a87cd",
  1026 => x"87d987c9",
  1027 => x"dbfa4973",
  1028 => x"7487d287",
  1029 => x"c149c01e",
  1030 => x"7487c7db",
  1031 => x"c149731e",
  1032 => x"c887ffda",
  1033 => x"87fbfd86",
  1034 => x"5c5b5e0e",
  1035 => x"711e0e5d",
  1036 => x"91de494c",
  1037 => x"4dfcecc2",
  1038 => x"6d978571",
  1039 => x"87dcc102",
  1040 => x"bfe8ecc2",
  1041 => x"7282744a",
  1042 => x"87ddfd49",
  1043 => x"026e7e70",
  1044 => x"c287f2c0",
  1045 => x"6e4bf0ec",
  1046 => x"ff49cb4a",
  1047 => x"7487c9c1",
  1048 => x"c193cb4b",
  1049 => x"c483cae3",
  1050 => x"e0c2c183",
  1051 => x"c149747b",
  1052 => x"7587ffc4",
  1053 => x"fbe2c17b",
  1054 => x"1e49bf97",
  1055 => x"49f0ecc2",
  1056 => x"c487e5fd",
  1057 => x"c1497486",
  1058 => x"c087e7c4",
  1059 => x"c6c6c149",
  1060 => x"d0ecc287",
  1061 => x"c178c048",
  1062 => x"87ffdc49",
  1063 => x"87c1fc26",
  1064 => x"64616f4c",
  1065 => x"2e676e69",
  1066 => x"0e002e2e",
  1067 => x"0e5c5b5e",
  1068 => x"c24a4b71",
  1069 => x"82bfe8ec",
  1070 => x"ecfb4972",
  1071 => x"9c4c7087",
  1072 => x"4987c402",
  1073 => x"c287dee7",
  1074 => x"c048e8ec",
  1075 => x"dc49c178",
  1076 => x"cefb87c9",
  1077 => x"5b5e0e87",
  1078 => x"f40e5d5c",
  1079 => x"dedfc286",
  1080 => x"c44cc04d",
  1081 => x"78c048a6",
  1082 => x"bfe8ecc2",
  1083 => x"06a9c049",
  1084 => x"c287c1c1",
  1085 => x"9848dedf",
  1086 => x"87f8c002",
  1087 => x"1efef7c0",
  1088 => x"c70266c8",
  1089 => x"48a6c487",
  1090 => x"87c578c0",
  1091 => x"c148a6c4",
  1092 => x"4966c478",
  1093 => x"c487c6e7",
  1094 => x"c14d7086",
  1095 => x"4866c484",
  1096 => x"a6c880c1",
  1097 => x"e8ecc258",
  1098 => x"03ac49bf",
  1099 => x"9d7587c6",
  1100 => x"87c8ff05",
  1101 => x"9d754cc0",
  1102 => x"87e0c302",
  1103 => x"1efef7c0",
  1104 => x"c70266c8",
  1105 => x"48a6cc87",
  1106 => x"87c578c0",
  1107 => x"c148a6cc",
  1108 => x"4966cc78",
  1109 => x"c487c6e6",
  1110 => x"6e7e7086",
  1111 => x"87e9c202",
  1112 => x"81cb496e",
  1113 => x"d0496997",
  1114 => x"d6c10299",
  1115 => x"ebc2c187",
  1116 => x"cb49744a",
  1117 => x"cae3c191",
  1118 => x"c8797281",
  1119 => x"51ffc381",
  1120 => x"91de4974",
  1121 => x"4dfcecc2",
  1122 => x"c1c28571",
  1123 => x"a5c17d97",
  1124 => x"51e0c049",
  1125 => x"97eee7c2",
  1126 => x"87d202bf",
  1127 => x"a5c284c1",
  1128 => x"eee7c24b",
  1129 => x"fe49db4a",
  1130 => x"c187fdfb",
  1131 => x"a5cd87db",
  1132 => x"c151c049",
  1133 => x"4ba5c284",
  1134 => x"49cb4a6e",
  1135 => x"87e8fbfe",
  1136 => x"c187c6c1",
  1137 => x"744ae8c0",
  1138 => x"c191cb49",
  1139 => x"7281cae3",
  1140 => x"eee7c279",
  1141 => x"d802bf97",
  1142 => x"de497487",
  1143 => x"c284c191",
  1144 => x"714bfcec",
  1145 => x"eee7c283",
  1146 => x"fe49dd4a",
  1147 => x"d887f9fa",
  1148 => x"de4b7487",
  1149 => x"fcecc293",
  1150 => x"49a3cb83",
  1151 => x"84c151c0",
  1152 => x"cb4a6e73",
  1153 => x"dffafe49",
  1154 => x"4866c487",
  1155 => x"a6c880c1",
  1156 => x"03acc758",
  1157 => x"6e87c5c0",
  1158 => x"87e0fc05",
  1159 => x"8ef44874",
  1160 => x"1e87fef5",
  1161 => x"4b711e73",
  1162 => x"c191cb49",
  1163 => x"c881cae3",
  1164 => x"e2c14aa1",
  1165 => x"501248fa",
  1166 => x"c04aa1c9",
  1167 => x"1248ebfa",
  1168 => x"c181ca50",
  1169 => x"1148fbe2",
  1170 => x"fbe2c150",
  1171 => x"1e49bf97",
  1172 => x"d3f649c0",
  1173 => x"d0ecc287",
  1174 => x"c178de48",
  1175 => x"87fbd549",
  1176 => x"87c1f526",
  1177 => x"494a711e",
  1178 => x"e3c191cb",
  1179 => x"81c881ca",
  1180 => x"ecc24811",
  1181 => x"ecc258d4",
  1182 => x"78c048e8",
  1183 => x"dad549c1",
  1184 => x"1e4f2687",
  1185 => x"fec049c0",
  1186 => x"4f2687cd",
  1187 => x"0299711e",
  1188 => x"e4c187d2",
  1189 => x"50c048df",
  1190 => x"c9c180f7",
  1191 => x"e3c140e4",
  1192 => x"87ce78c3",
  1193 => x"48dbe4c1",
  1194 => x"78fce2c1",
  1195 => x"cac180fc",
  1196 => x"4f2678c3",
  1197 => x"5c5b5e0e",
  1198 => x"4a4c710e",
  1199 => x"e3c192cb",
  1200 => x"a2c882ca",
  1201 => x"4ba2c949",
  1202 => x"1e4b6b97",
  1203 => x"1e496997",
  1204 => x"491282ca",
  1205 => x"87c6e7c0",
  1206 => x"fed349c0",
  1207 => x"c0497487",
  1208 => x"f887cffb",
  1209 => x"87fbf28e",
  1210 => x"711e731e",
  1211 => x"c3ff494b",
  1212 => x"fe497387",
  1213 => x"ecf287fe",
  1214 => x"1e731e87",
  1215 => x"a3c64b71",
  1216 => x"87db024a",
  1217 => x"d6028ac1",
  1218 => x"c1028a87",
  1219 => x"028a87da",
  1220 => x"8a87fcc0",
  1221 => x"87e1c002",
  1222 => x"87cb028a",
  1223 => x"c787dbc1",
  1224 => x"87c0fd49",
  1225 => x"c287dec1",
  1226 => x"02bfe8ec",
  1227 => x"4887cbc1",
  1228 => x"ecc288c1",
  1229 => x"c1c158ec",
  1230 => x"ececc287",
  1231 => x"f9c002bf",
  1232 => x"e8ecc287",
  1233 => x"80c148bf",
  1234 => x"58ececc2",
  1235 => x"c287ebc0",
  1236 => x"49bfe8ec",
  1237 => x"ecc289c6",
  1238 => x"b7c059ec",
  1239 => x"87da03a9",
  1240 => x"48e8ecc2",
  1241 => x"87d278c0",
  1242 => x"bfececc2",
  1243 => x"c287cb02",
  1244 => x"48bfe8ec",
  1245 => x"ecc280c6",
  1246 => x"49c058ec",
  1247 => x"7387dcd1",
  1248 => x"edf8c049",
  1249 => x"87ddf087",
  1250 => x"5c5b5e0e",
  1251 => x"cc4c710e",
  1252 => x"4b741e66",
  1253 => x"e3c193cb",
  1254 => x"a3c483ca",
  1255 => x"fe496a4a",
  1256 => x"c187d5f4",
  1257 => x"c87be3c8",
  1258 => x"66d449a3",
  1259 => x"49a3c951",
  1260 => x"ca5166d8",
  1261 => x"66dc49a3",
  1262 => x"e6ef2651",
  1263 => x"5b5e0e87",
  1264 => x"ff0e5d5c",
  1265 => x"a6d886d0",
  1266 => x"48a6c459",
  1267 => x"80c478c0",
  1268 => x"7866c4c1",
  1269 => x"78c180c4",
  1270 => x"78c180c4",
  1271 => x"48ececc2",
  1272 => x"ecc278c1",
  1273 => x"de48bfd0",
  1274 => x"87cb05a8",
  1275 => x"7087e6f3",
  1276 => x"59a6c849",
  1277 => x"e387ecce",
  1278 => x"c9e487e7",
  1279 => x"87d6e387",
  1280 => x"fbc04c70",
  1281 => x"d0c102ac",
  1282 => x"0566d487",
  1283 => x"c087c2c1",
  1284 => x"1ec11e1e",
  1285 => x"1efde4c1",
  1286 => x"ebfd49c0",
  1287 => x"66d0c187",
  1288 => x"6a82c44a",
  1289 => x"7481c749",
  1290 => x"d81ec151",
  1291 => x"c8496a1e",
  1292 => x"87e6e381",
  1293 => x"c4c186d8",
  1294 => x"a8c04866",
  1295 => x"c487c701",
  1296 => x"78c148a6",
  1297 => x"c4c187ce",
  1298 => x"88c14866",
  1299 => x"c358a6cc",
  1300 => x"87f2e287",
  1301 => x"c248a6cc",
  1302 => x"029c7478",
  1303 => x"c487c0cd",
  1304 => x"c8c14866",
  1305 => x"cc03a866",
  1306 => x"a6d887f5",
  1307 => x"c478c048",
  1308 => x"e178c080",
  1309 => x"4c7087e0",
  1310 => x"05acd0c1",
  1311 => x"dc87d8c2",
  1312 => x"c4e47e66",
  1313 => x"c0497087",
  1314 => x"e159a6e0",
  1315 => x"4c7087c8",
  1316 => x"05acecc0",
  1317 => x"c487ebc1",
  1318 => x"91cb4966",
  1319 => x"8166c0c1",
  1320 => x"6a4aa1c4",
  1321 => x"4aa1c84d",
  1322 => x"c15266dc",
  1323 => x"e079e4c9",
  1324 => x"4c7087e4",
  1325 => x"87d8029c",
  1326 => x"02acfbc0",
  1327 => x"557487d2",
  1328 => x"7087d3e0",
  1329 => x"c7029c4c",
  1330 => x"acfbc087",
  1331 => x"87eeff05",
  1332 => x"c255e0c0",
  1333 => x"97c055c1",
  1334 => x"4966d47d",
  1335 => x"db05a96e",
  1336 => x"4866c487",
  1337 => x"04a866c8",
  1338 => x"66c487ca",
  1339 => x"c880c148",
  1340 => x"87c858a6",
  1341 => x"c14866c8",
  1342 => x"58a6cc88",
  1343 => x"87d6dfff",
  1344 => x"d0c14c70",
  1345 => x"87c805ac",
  1346 => x"c14866d0",
  1347 => x"58a6d480",
  1348 => x"02acd0c1",
  1349 => x"c087e8fd",
  1350 => x"d448a6e0",
  1351 => x"66dc7866",
  1352 => x"66e0c048",
  1353 => x"c8c905a8",
  1354 => x"a6e4c087",
  1355 => x"7e78c048",
  1356 => x"fbc04874",
  1357 => x"a6ecc088",
  1358 => x"02987058",
  1359 => x"4887cdc8",
  1360 => x"ecc088cb",
  1361 => x"987058a6",
  1362 => x"87d2c102",
  1363 => x"c088c948",
  1364 => x"7058a6ec",
  1365 => x"dbc30298",
  1366 => x"88c44887",
  1367 => x"58a6ecc0",
  1368 => x"d0029870",
  1369 => x"88c14887",
  1370 => x"58a6ecc0",
  1371 => x"c3029870",
  1372 => x"d1c787c2",
  1373 => x"48a6d887",
  1374 => x"ff78f0c0",
  1375 => x"7087d7dd",
  1376 => x"acecc04c",
  1377 => x"87c3c002",
  1378 => x"c05ca6dc",
  1379 => x"cd02acec",
  1380 => x"c1ddff87",
  1381 => x"c04c7087",
  1382 => x"ff05acec",
  1383 => x"ecc087f3",
  1384 => x"c4c002ac",
  1385 => x"eddcff87",
  1386 => x"1e66d887",
  1387 => x"1e4966d4",
  1388 => x"1e4966d4",
  1389 => x"1efde4c1",
  1390 => x"f74966d4",
  1391 => x"1ec087ca",
  1392 => x"66dc1eca",
  1393 => x"c191cb49",
  1394 => x"d88166d8",
  1395 => x"a1c448a6",
  1396 => x"bf66d878",
  1397 => x"c1ddff49",
  1398 => x"c086d887",
  1399 => x"c106a8b7",
  1400 => x"1ec187c5",
  1401 => x"66c81ede",
  1402 => x"dcff49bf",
  1403 => x"86c887ec",
  1404 => x"c0484970",
  1405 => x"a6dc8808",
  1406 => x"a8b7c058",
  1407 => x"87e7c006",
  1408 => x"dd4866d8",
  1409 => x"de03a8b7",
  1410 => x"49bf6e87",
  1411 => x"c08166d8",
  1412 => x"66d851e0",
  1413 => x"6e81c149",
  1414 => x"c1c281bf",
  1415 => x"4966d851",
  1416 => x"bf6e81c2",
  1417 => x"cc51c081",
  1418 => x"80c14866",
  1419 => x"c158a6d0",
  1420 => x"87d8c47e",
  1421 => x"87d1ddff",
  1422 => x"ff58a6dc",
  1423 => x"c087cadd",
  1424 => x"c058a6ec",
  1425 => x"c005a8ec",
  1426 => x"e8c087ca",
  1427 => x"66d848a6",
  1428 => x"87c4c078",
  1429 => x"87fed9ff",
  1430 => x"cb4966c4",
  1431 => x"66c0c191",
  1432 => x"70807148",
  1433 => x"c8496e7e",
  1434 => x"ca4a6e81",
  1435 => x"5266d882",
  1436 => x"4a66e8c0",
  1437 => x"66d882c1",
  1438 => x"7248c18a",
  1439 => x"c14a7030",
  1440 => x"7997728a",
  1441 => x"1e496997",
  1442 => x"d74966dc",
  1443 => x"86c487d2",
  1444 => x"58a6f0c0",
  1445 => x"81c4496e",
  1446 => x"e0c04d69",
  1447 => x"66dc4866",
  1448 => x"c8c002a8",
  1449 => x"48a6d887",
  1450 => x"c5c078c0",
  1451 => x"48a6d887",
  1452 => x"66d878c1",
  1453 => x"1ee0c01e",
  1454 => x"d9ff4975",
  1455 => x"86c887dc",
  1456 => x"b7c04c70",
  1457 => x"d4c106ac",
  1458 => x"c0857487",
  1459 => x"897449e0",
  1460 => x"dfc14b75",
  1461 => x"fe714ad8",
  1462 => x"c287cde7",
  1463 => x"66e4c085",
  1464 => x"c080c148",
  1465 => x"c058a6e8",
  1466 => x"c14966ec",
  1467 => x"02a97081",
  1468 => x"d887c8c0",
  1469 => x"78c048a6",
  1470 => x"d887c5c0",
  1471 => x"78c148a6",
  1472 => x"c21e66d8",
  1473 => x"e0c049a4",
  1474 => x"70887148",
  1475 => x"49751e49",
  1476 => x"87c6d8ff",
  1477 => x"b7c086c8",
  1478 => x"c0ff01a8",
  1479 => x"66e4c087",
  1480 => x"87d1c002",
  1481 => x"81c9496e",
  1482 => x"5166e4c0",
  1483 => x"cac1486e",
  1484 => x"ccc078f4",
  1485 => x"c9496e87",
  1486 => x"6e51c281",
  1487 => x"e8cbc148",
  1488 => x"c07ec178",
  1489 => x"d6ff87c6",
  1490 => x"4c7087fc",
  1491 => x"f5c0026e",
  1492 => x"4866c487",
  1493 => x"04a866c8",
  1494 => x"c487cbc0",
  1495 => x"80c14866",
  1496 => x"c058a6c8",
  1497 => x"66c887e0",
  1498 => x"cc88c148",
  1499 => x"d5c058a6",
  1500 => x"acc6c187",
  1501 => x"87c8c005",
  1502 => x"c14866cc",
  1503 => x"58a6d080",
  1504 => x"87c2d6ff",
  1505 => x"66d04c70",
  1506 => x"d480c148",
  1507 => x"9c7458a6",
  1508 => x"87cbc002",
  1509 => x"c14866c4",
  1510 => x"04a866c8",
  1511 => x"ff87cbf3",
  1512 => x"c487dad5",
  1513 => x"a8c74866",
  1514 => x"87e5c003",
  1515 => x"48ececc2",
  1516 => x"66c478c0",
  1517 => x"c191cb49",
  1518 => x"c48166c0",
  1519 => x"4a6a4aa1",
  1520 => x"c47952c0",
  1521 => x"80c14866",
  1522 => x"c758a6c8",
  1523 => x"dbff04a8",
  1524 => x"8ed0ff87",
  1525 => x"87c9dfff",
  1526 => x"1e00203a",
  1527 => x"4b711e73",
  1528 => x"87c6029b",
  1529 => x"48e8ecc2",
  1530 => x"1ec778c0",
  1531 => x"bfe8ecc2",
  1532 => x"e3c11e49",
  1533 => x"ecc21eca",
  1534 => x"ee49bfd0",
  1535 => x"86cc87ff",
  1536 => x"bfd0ecc2",
  1537 => x"87c4ea49",
  1538 => x"c8029b73",
  1539 => x"cae3c187",
  1540 => x"efe7c049",
  1541 => x"ccdeff87",
  1542 => x"e2c11e87",
  1543 => x"50c048fa",
  1544 => x"bfede4c1",
  1545 => x"c3daff49",
  1546 => x"2648c087",
  1547 => x"ebc71e4f",
  1548 => x"fe49c187",
  1549 => x"eafe87e5",
  1550 => x"987087e3",
  1551 => x"fe87cd02",
  1552 => x"7087def3",
  1553 => x"87c40298",
  1554 => x"87c24ac1",
  1555 => x"9a724ac0",
  1556 => x"c087ce05",
  1557 => x"c1e2c11e",
  1558 => x"fff2c049",
  1559 => x"fe86c487",
  1560 => x"e7fcc087",
  1561 => x"c11ec087",
  1562 => x"c049cce2",
  1563 => x"c087edf2",
  1564 => x"87e5fe1e",
  1565 => x"f2c04970",
  1566 => x"dec387e2",
  1567 => x"268ef887",
  1568 => x"2044534f",
  1569 => x"6c696166",
  1570 => x"002e6465",
  1571 => x"746f6f42",
  1572 => x"2e676e69",
  1573 => x"1e002e2e",
  1574 => x"87c4eac0",
  1575 => x"87f2f5c0",
  1576 => x"4f2687f6",
  1577 => x"e8ecc21e",
  1578 => x"c278c048",
  1579 => x"c048d0ec",
  1580 => x"87f9fd78",
  1581 => x"48c087e1",
  1582 => x"00004f26",
  1583 => x"78452080",
  1584 => x"80007469",
  1585 => x"63614220",
  1586 => x"1264006b",
  1587 => x"2b3c0000",
  1588 => x"00000000",
  1589 => x"00126400",
  1590 => x"002b5a00",
  1591 => x"00000000",
  1592 => x"00001264",
  1593 => x"00002b78",
  1594 => x"64000000",
  1595 => x"96000012",
  1596 => x"0000002b",
  1597 => x"12640000",
  1598 => x"2bb40000",
  1599 => x"00000000",
  1600 => x"00126400",
  1601 => x"002bd200",
  1602 => x"00000000",
  1603 => x"00001264",
  1604 => x"00002bf0",
  1605 => x"64000000",
  1606 => x"00000012",
  1607 => x"00000000",
  1608 => x"12f90000",
  1609 => x"00000000",
  1610 => x"00000000",
  1611 => x"00193100",
  1612 => x"34364300",
  1613 => x"20202020",
  1614 => x"4d4f5220",
  1615 => x"616f4c00",
  1616 => x"2e2a2064",
  1617 => x"f0fe1e00",
  1618 => x"cd78c048",
  1619 => x"26097909",
  1620 => x"fe1e1e4f",
  1621 => x"487ebff0",
  1622 => x"1e4f2626",
  1623 => x"c148f0fe",
  1624 => x"1e4f2678",
  1625 => x"c048f0fe",
  1626 => x"1e4f2678",
  1627 => x"52c04a71",
  1628 => x"0e4f2652",
  1629 => x"5d5c5b5e",
  1630 => x"7186f40e",
  1631 => x"7e6d974d",
  1632 => x"974ca5c1",
  1633 => x"a6c8486c",
  1634 => x"c4486e58",
  1635 => x"c505a866",
  1636 => x"c048ff87",
  1637 => x"caff87e6",
  1638 => x"49a5c287",
  1639 => x"714b6c97",
  1640 => x"6b974ba3",
  1641 => x"7e6c974b",
  1642 => x"80c1486e",
  1643 => x"c758a6c8",
  1644 => x"58a6cc98",
  1645 => x"fe7c9770",
  1646 => x"487387e1",
  1647 => x"4d268ef4",
  1648 => x"4b264c26",
  1649 => x"5e0e4f26",
  1650 => x"f40e5c5b",
  1651 => x"d84c7186",
  1652 => x"ffc34a66",
  1653 => x"4ba4c29a",
  1654 => x"73496c97",
  1655 => x"517249a1",
  1656 => x"6e7e6c97",
  1657 => x"c880c148",
  1658 => x"98c758a6",
  1659 => x"7058a6cc",
  1660 => x"ff8ef454",
  1661 => x"1e1e87ca",
  1662 => x"e087e8fd",
  1663 => x"c0494abf",
  1664 => x"0299c0e0",
  1665 => x"1e7287cb",
  1666 => x"49cef0c2",
  1667 => x"c487f7fe",
  1668 => x"87fdfc86",
  1669 => x"c2fd7e70",
  1670 => x"4f262687",
  1671 => x"cef0c21e",
  1672 => x"87c7fd49",
  1673 => x"49f6e7c1",
  1674 => x"c487dafc",
  1675 => x"4f2687c7",
  1676 => x"48d0ff1e",
  1677 => x"ff78e1c8",
  1678 => x"78c548d4",
  1679 => x"c30266c4",
  1680 => x"78e0c387",
  1681 => x"c60266c8",
  1682 => x"48d4ff87",
  1683 => x"ff78f0c3",
  1684 => x"787148d4",
  1685 => x"c848d0ff",
  1686 => x"e0c078e1",
  1687 => x"0e4f2678",
  1688 => x"0e5c5b5e",
  1689 => x"f0c24c71",
  1690 => x"c6fc49ce",
  1691 => x"c04a7087",
  1692 => x"c204aab7",
  1693 => x"f0c387e2",
  1694 => x"87c905aa",
  1695 => x"48e4ecc1",
  1696 => x"c3c278c1",
  1697 => x"aae0c387",
  1698 => x"c187c905",
  1699 => x"c148e8ec",
  1700 => x"87f4c178",
  1701 => x"bfe8ecc1",
  1702 => x"c287c602",
  1703 => x"c24ba2c0",
  1704 => x"744b7287",
  1705 => x"87d1059c",
  1706 => x"bfe4ecc1",
  1707 => x"e8ecc11e",
  1708 => x"49721ebf",
  1709 => x"c887f9fd",
  1710 => x"e4ecc186",
  1711 => x"e0c002bf",
  1712 => x"c4497387",
  1713 => x"c19129b7",
  1714 => x"7381c4ee",
  1715 => x"c29acf4a",
  1716 => x"7248c192",
  1717 => x"ff4a7030",
  1718 => x"694872ba",
  1719 => x"db797098",
  1720 => x"c4497387",
  1721 => x"c19129b7",
  1722 => x"7381c4ee",
  1723 => x"c29acf4a",
  1724 => x"7248c392",
  1725 => x"484a7030",
  1726 => x"7970b069",
  1727 => x"48e8ecc1",
  1728 => x"ecc178c0",
  1729 => x"78c048e4",
  1730 => x"49cef0c2",
  1731 => x"7087e4f9",
  1732 => x"aab7c04a",
  1733 => x"87defd03",
  1734 => x"87c248c0",
  1735 => x"4c264d26",
  1736 => x"4f264b26",
  1737 => x"00000000",
  1738 => x"00000000",
  1739 => x"494a711e",
  1740 => x"2687ecfc",
  1741 => x"4ac01e4f",
  1742 => x"91c44972",
  1743 => x"81c4eec1",
  1744 => x"82c179c0",
  1745 => x"04aab7d0",
  1746 => x"4f2687ee",
  1747 => x"5c5b5e0e",
  1748 => x"4d710e5d",
  1749 => x"7587ccf8",
  1750 => x"2ab7c44a",
  1751 => x"c4eec192",
  1752 => x"cf4c7582",
  1753 => x"6a94c29c",
  1754 => x"2b744b49",
  1755 => x"48c29bc3",
  1756 => x"4c703074",
  1757 => x"4874bcff",
  1758 => x"7a709871",
  1759 => x"7387dcf7",
  1760 => x"87d8fe48",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"48d0ff1e",
  1778 => x"7178e1c8",
  1779 => x"08d4ff48",
  1780 => x"1e4f2678",
  1781 => x"c848d0ff",
  1782 => x"487178e1",
  1783 => x"7808d4ff",
  1784 => x"ff4866c4",
  1785 => x"267808d4",
  1786 => x"4a711e4f",
  1787 => x"1e4966c4",
  1788 => x"deff4972",
  1789 => x"48d0ff87",
  1790 => x"2678e0c0",
  1791 => x"731e4f26",
  1792 => x"c84b711e",
  1793 => x"731e4966",
  1794 => x"a2e0c14a",
  1795 => x"87d9ff49",
  1796 => x"2687c426",
  1797 => x"264c264d",
  1798 => x"1e4f264b",
  1799 => x"c34ad4ff",
  1800 => x"d0ff7aff",
  1801 => x"78e1c048",
  1802 => x"f0c27ade",
  1803 => x"497abfd8",
  1804 => x"7028c848",
  1805 => x"d048717a",
  1806 => x"717a7028",
  1807 => x"7028d848",
  1808 => x"dcf0c27a",
  1809 => x"48497abf",
  1810 => x"7a7028c8",
  1811 => x"28d04871",
  1812 => x"48717a70",
  1813 => x"7a7028d8",
  1814 => x"c048d0ff",
  1815 => x"4f2678e0",
  1816 => x"711e731e",
  1817 => x"d8f0c24a",
  1818 => x"2b724bbf",
  1819 => x"04aae0c0",
  1820 => x"497287ce",
  1821 => x"c289e0c0",
  1822 => x"4bbfdcf0",
  1823 => x"87cf2b71",
  1824 => x"7249e0c0",
  1825 => x"dcf0c289",
  1826 => x"307148bf",
  1827 => x"c8b34970",
  1828 => x"48739b66",
  1829 => x"4d2687c4",
  1830 => x"4b264c26",
  1831 => x"5e0e4f26",
  1832 => x"0e5d5c5b",
  1833 => x"4b7186ec",
  1834 => x"bfd8f0c2",
  1835 => x"2c734c7e",
  1836 => x"04abe0c0",
  1837 => x"c487e0c0",
  1838 => x"78c048a6",
  1839 => x"e0c04973",
  1840 => x"c04a7189",
  1841 => x"724866e4",
  1842 => x"58a6cc30",
  1843 => x"bfdcf0c2",
  1844 => x"2c714c4d",
  1845 => x"7387e4c0",
  1846 => x"66e4c049",
  1847 => x"c8307148",
  1848 => x"e0c058a6",
  1849 => x"c0897349",
  1850 => x"714866e4",
  1851 => x"58a6cc28",
  1852 => x"bfdcf0c2",
  1853 => x"3071484d",
  1854 => x"c0b44970",
  1855 => x"c19c66e4",
  1856 => x"66e8c084",
  1857 => x"87c204ac",
  1858 => x"e0c04cc0",
  1859 => x"87d304ab",
  1860 => x"c048a6cc",
  1861 => x"c0497378",
  1862 => x"487489e0",
  1863 => x"a6d43071",
  1864 => x"7387d558",
  1865 => x"71487449",
  1866 => x"58a6d030",
  1867 => x"7349e0c0",
  1868 => x"71487489",
  1869 => x"58a6d428",
  1870 => x"ff4a66c4",
  1871 => x"c89a6eba",
  1872 => x"b9ff4966",
  1873 => x"48729975",
  1874 => x"c2b066cc",
  1875 => x"7158dcf0",
  1876 => x"b066d048",
  1877 => x"58e0f0c2",
  1878 => x"ec87c0fb",
  1879 => x"87f6fc8e",
  1880 => x"48d0ff1e",
  1881 => x"7178c9c8",
  1882 => x"08d4ff48",
  1883 => x"1e4f2678",
  1884 => x"eb494a71",
  1885 => x"48d0ff87",
  1886 => x"4f2678c8",
  1887 => x"711e731e",
  1888 => x"ecf0c24b",
  1889 => x"87c302bf",
  1890 => x"ff87ebc2",
  1891 => x"c9c848d0",
  1892 => x"c0497378",
  1893 => x"d4ffb1e0",
  1894 => x"c2787148",
  1895 => x"c048e0f0",
  1896 => x"0266c878",
  1897 => x"ffc387c5",
  1898 => x"c087c249",
  1899 => x"e8f0c249",
  1900 => x"0266cc59",
  1901 => x"d5c587c6",
  1902 => x"87c44ad5",
  1903 => x"4affffcf",
  1904 => x"5aecf0c2",
  1905 => x"48ecf0c2",
  1906 => x"87c478c1",
  1907 => x"4c264d26",
  1908 => x"4f264b26",
  1909 => x"5c5b5e0e",
  1910 => x"4a710e5d",
  1911 => x"bfe8f0c2",
  1912 => x"029a724c",
  1913 => x"c84987cb",
  1914 => x"f2f5c191",
  1915 => x"c483714b",
  1916 => x"f2f9c187",
  1917 => x"134dc04b",
  1918 => x"c2997449",
  1919 => x"b9bfe4f0",
  1920 => x"7148d4ff",
  1921 => x"2cb7c178",
  1922 => x"adb7c885",
  1923 => x"c287e804",
  1924 => x"48bfe0f0",
  1925 => x"f0c280c8",
  1926 => x"effe58e4",
  1927 => x"1e731e87",
  1928 => x"4a134b71",
  1929 => x"87cb029a",
  1930 => x"e7fe4972",
  1931 => x"9a4a1387",
  1932 => x"fe87f505",
  1933 => x"c21e87da",
  1934 => x"49bfe0f0",
  1935 => x"48e0f0c2",
  1936 => x"c478a1c1",
  1937 => x"03a9b7c0",
  1938 => x"d4ff87db",
  1939 => x"e4f0c248",
  1940 => x"f0c278bf",
  1941 => x"c249bfe0",
  1942 => x"c148e0f0",
  1943 => x"c0c478a1",
  1944 => x"e504a9b7",
  1945 => x"48d0ff87",
  1946 => x"f0c278c8",
  1947 => x"78c048ec",
  1948 => x"00004f26",
  1949 => x"00000000",
  1950 => x"00000000",
  1951 => x"005f5f00",
  1952 => x"03000000",
  1953 => x"03030003",
  1954 => x"7f140000",
  1955 => x"7f7f147f",
  1956 => x"24000014",
  1957 => x"3a6b6b2e",
  1958 => x"6a4c0012",
  1959 => x"566c1836",
  1960 => x"7e300032",
  1961 => x"3a77594f",
  1962 => x"00004068",
  1963 => x"00030704",
  1964 => x"00000000",
  1965 => x"41633e1c",
  1966 => x"00000000",
  1967 => x"1c3e6341",
  1968 => x"2a080000",
  1969 => x"3e1c1c3e",
  1970 => x"0800082a",
  1971 => x"083e3e08",
  1972 => x"00000008",
  1973 => x"0060e080",
  1974 => x"08000000",
  1975 => x"08080808",
  1976 => x"00000008",
  1977 => x"00606000",
  1978 => x"60400000",
  1979 => x"060c1830",
  1980 => x"3e000103",
  1981 => x"7f4d597f",
  1982 => x"0400003e",
  1983 => x"007f7f06",
  1984 => x"42000000",
  1985 => x"4f597163",
  1986 => x"22000046",
  1987 => x"7f494963",
  1988 => x"1c180036",
  1989 => x"7f7f1316",
  1990 => x"27000010",
  1991 => x"7d454567",
  1992 => x"3c000039",
  1993 => x"79494b7e",
  1994 => x"01000030",
  1995 => x"0f797101",
  1996 => x"36000007",
  1997 => x"7f49497f",
  1998 => x"06000036",
  1999 => x"3f69494f",
  2000 => x"0000001e",
  2001 => x"00666600",
  2002 => x"00000000",
  2003 => x"0066e680",
  2004 => x"08000000",
  2005 => x"22141408",
  2006 => x"14000022",
  2007 => x"14141414",
  2008 => x"22000014",
  2009 => x"08141422",
  2010 => x"02000008",
  2011 => x"0f595103",
  2012 => x"7f3e0006",
  2013 => x"1f555d41",
  2014 => x"7e00001e",
  2015 => x"7f09097f",
  2016 => x"7f00007e",
  2017 => x"7f49497f",
  2018 => x"1c000036",
  2019 => x"4141633e",
  2020 => x"7f000041",
  2021 => x"3e63417f",
  2022 => x"7f00001c",
  2023 => x"4149497f",
  2024 => x"7f000041",
  2025 => x"0109097f",
  2026 => x"3e000001",
  2027 => x"7b49417f",
  2028 => x"7f00007a",
  2029 => x"7f08087f",
  2030 => x"0000007f",
  2031 => x"417f7f41",
  2032 => x"20000000",
  2033 => x"7f404060",
  2034 => x"7f7f003f",
  2035 => x"63361c08",
  2036 => x"7f000041",
  2037 => x"4040407f",
  2038 => x"7f7f0040",
  2039 => x"7f060c06",
  2040 => x"7f7f007f",
  2041 => x"7f180c06",
  2042 => x"3e00007f",
  2043 => x"7f41417f",
  2044 => x"7f00003e",
  2045 => x"0f09097f",
  2046 => x"7f3e0006",
  2047 => x"7e7f6141",
  2048 => x"7f000040",
  2049 => x"7f19097f",
  2050 => x"26000066",
  2051 => x"7b594d6f",
  2052 => x"01000032",
  2053 => x"017f7f01",
  2054 => x"3f000001",
  2055 => x"7f40407f",
  2056 => x"0f00003f",
  2057 => x"3f70703f",
  2058 => x"7f7f000f",
  2059 => x"7f301830",
  2060 => x"6341007f",
  2061 => x"361c1c36",
  2062 => x"03014163",
  2063 => x"067c7c06",
  2064 => x"71610103",
  2065 => x"43474d59",
  2066 => x"00000041",
  2067 => x"41417f7f",
  2068 => x"03010000",
  2069 => x"30180c06",
  2070 => x"00004060",
  2071 => x"7f7f4141",
  2072 => x"0c080000",
  2073 => x"0c060306",
  2074 => x"80800008",
  2075 => x"80808080",
  2076 => x"00000080",
  2077 => x"04070300",
  2078 => x"20000000",
  2079 => x"7c545474",
  2080 => x"7f000078",
  2081 => x"7c44447f",
  2082 => x"38000038",
  2083 => x"4444447c",
  2084 => x"38000000",
  2085 => x"7f44447c",
  2086 => x"3800007f",
  2087 => x"5c54547c",
  2088 => x"04000018",
  2089 => x"05057f7e",
  2090 => x"18000000",
  2091 => x"fca4a4bc",
  2092 => x"7f00007c",
  2093 => x"7c04047f",
  2094 => x"00000078",
  2095 => x"407d3d00",
  2096 => x"80000000",
  2097 => x"7dfd8080",
  2098 => x"7f000000",
  2099 => x"6c38107f",
  2100 => x"00000044",
  2101 => x"407f3f00",
  2102 => x"7c7c0000",
  2103 => x"7c0c180c",
  2104 => x"7c000078",
  2105 => x"7c04047c",
  2106 => x"38000078",
  2107 => x"7c44447c",
  2108 => x"fc000038",
  2109 => x"3c2424fc",
  2110 => x"18000018",
  2111 => x"fc24243c",
  2112 => x"7c0000fc",
  2113 => x"0c04047c",
  2114 => x"48000008",
  2115 => x"7454545c",
  2116 => x"04000020",
  2117 => x"44447f3f",
  2118 => x"3c000000",
  2119 => x"7c40407c",
  2120 => x"1c00007c",
  2121 => x"3c60603c",
  2122 => x"7c3c001c",
  2123 => x"7c603060",
  2124 => x"6c44003c",
  2125 => x"6c381038",
  2126 => x"1c000044",
  2127 => x"3c60e0bc",
  2128 => x"4400001c",
  2129 => x"4c5c7464",
  2130 => x"08000044",
  2131 => x"41773e08",
  2132 => x"00000041",
  2133 => x"007f7f00",
  2134 => x"41000000",
  2135 => x"083e7741",
  2136 => x"01020008",
  2137 => x"02020301",
  2138 => x"7f7f0001",
  2139 => x"7f7f7f7f",
  2140 => x"0808007f",
  2141 => x"3e3e1c1c",
  2142 => x"7f7f7f7f",
  2143 => x"1c1c3e3e",
  2144 => x"10000808",
  2145 => x"187c7c18",
  2146 => x"10000010",
  2147 => x"307c7c30",
  2148 => x"30100010",
  2149 => x"1e786060",
  2150 => x"66420006",
  2151 => x"663c183c",
  2152 => x"38780042",
  2153 => x"6cc6c26a",
  2154 => x"00600038",
  2155 => x"00006000",
  2156 => x"5e0e0060",
  2157 => x"0e5d5c5b",
  2158 => x"c24c711e",
  2159 => x"4dbffdf0",
  2160 => x"1ec04bc0",
  2161 => x"c702ab74",
  2162 => x"48a6c487",
  2163 => x"87c578c0",
  2164 => x"c148a6c4",
  2165 => x"1e66c478",
  2166 => x"dfee4973",
  2167 => x"c086c887",
  2168 => x"efef49e0",
  2169 => x"4aa5c487",
  2170 => x"f0f0496a",
  2171 => x"87c6f187",
  2172 => x"83c185cb",
  2173 => x"04abb7c8",
  2174 => x"2687c7ff",
  2175 => x"4c264d26",
  2176 => x"4f264b26",
  2177 => x"c24a711e",
  2178 => x"c25ac1f1",
  2179 => x"c748c1f1",
  2180 => x"ddfe4978",
  2181 => x"1e4f2687",
  2182 => x"4a711e73",
  2183 => x"03aab7c0",
  2184 => x"d5c287d3",
  2185 => x"c405bff1",
  2186 => x"c24bc187",
  2187 => x"c24bc087",
  2188 => x"c45bf5d5",
  2189 => x"f5d5c287",
  2190 => x"f1d5c25a",
  2191 => x"9ac14abf",
  2192 => x"49a2c0c1",
  2193 => x"fc87e8ec",
  2194 => x"f1d5c248",
  2195 => x"effe78bf",
  2196 => x"4a711e87",
  2197 => x"721e66c4",
  2198 => x"87e2e649",
  2199 => x"1e4f2626",
  2200 => x"bff1d5c2",
  2201 => x"87c4e349",
  2202 => x"48f5f0c2",
  2203 => x"c278bfe8",
  2204 => x"ec48f1f0",
  2205 => x"f0c278bf",
  2206 => x"494abff5",
  2207 => x"c899ffc3",
  2208 => x"48722ab7",
  2209 => x"f0c2b071",
  2210 => x"4f2658fd",
  2211 => x"5c5b5e0e",
  2212 => x"4b710e5d",
  2213 => x"c287c8ff",
  2214 => x"c048f0f0",
  2215 => x"e2497350",
  2216 => x"497087ea",
  2217 => x"cb9cc24c",
  2218 => x"cccb49ee",
  2219 => x"4d497087",
  2220 => x"97f0f0c2",
  2221 => x"e2c105bf",
  2222 => x"4966d087",
  2223 => x"bff9f0c2",
  2224 => x"87d60599",
  2225 => x"c24966d4",
  2226 => x"99bff1f0",
  2227 => x"7387cb05",
  2228 => x"87f8e149",
  2229 => x"c1029870",
  2230 => x"4cc187c1",
  2231 => x"7587c0fe",
  2232 => x"87e1ca49",
  2233 => x"c6029870",
  2234 => x"f0f0c287",
  2235 => x"c250c148",
  2236 => x"bf97f0f0",
  2237 => x"87e3c005",
  2238 => x"bff9f0c2",
  2239 => x"9966d049",
  2240 => x"87d6ff05",
  2241 => x"bff1f0c2",
  2242 => x"9966d449",
  2243 => x"87caff05",
  2244 => x"f7e04973",
  2245 => x"05987087",
  2246 => x"7487fffe",
  2247 => x"87dcfb48",
  2248 => x"5c5b5e0e",
  2249 => x"86f40e5d",
  2250 => x"ec4c4dc0",
  2251 => x"a6c47ebf",
  2252 => x"fdf0c248",
  2253 => x"1ec178bf",
  2254 => x"49c71ec0",
  2255 => x"c887cdfd",
  2256 => x"02987086",
  2257 => x"49ff87ce",
  2258 => x"c187ccfb",
  2259 => x"dfff49da",
  2260 => x"4dc187fa",
  2261 => x"97f0f0c2",
  2262 => x"87c302bf",
  2263 => x"c287c4d0",
  2264 => x"4bbff5f0",
  2265 => x"bff1d5c2",
  2266 => x"87ebc005",
  2267 => x"ff49fdc3",
  2268 => x"c387d9df",
  2269 => x"dfff49fa",
  2270 => x"497387d2",
  2271 => x"7199ffc3",
  2272 => x"fb49c01e",
  2273 => x"497387cb",
  2274 => x"7129b7c8",
  2275 => x"fa49c11e",
  2276 => x"86c887ff",
  2277 => x"c287c0c6",
  2278 => x"4bbff9f0",
  2279 => x"87dd029b",
  2280 => x"bfedd5c2",
  2281 => x"87ddc749",
  2282 => x"c4059870",
  2283 => x"d24bc087",
  2284 => x"49e0c287",
  2285 => x"c287c2c7",
  2286 => x"c658f1d5",
  2287 => x"edd5c287",
  2288 => x"7378c048",
  2289 => x"0599c249",
  2290 => x"ebc387ce",
  2291 => x"fbddff49",
  2292 => x"c2497087",
  2293 => x"87c20299",
  2294 => x"49734cfb",
  2295 => x"ce0599c1",
  2296 => x"49f4c387",
  2297 => x"87e4ddff",
  2298 => x"99c24970",
  2299 => x"fa87c202",
  2300 => x"c849734c",
  2301 => x"87ce0599",
  2302 => x"ff49f5c3",
  2303 => x"7087cddd",
  2304 => x"0299c249",
  2305 => x"f1c287d5",
  2306 => x"ca02bfc1",
  2307 => x"88c14887",
  2308 => x"58c5f1c2",
  2309 => x"ff87c2c0",
  2310 => x"734dc14c",
  2311 => x"0599c449",
  2312 => x"f2c387ce",
  2313 => x"e3dcff49",
  2314 => x"c2497087",
  2315 => x"87dc0299",
  2316 => x"bfc1f1c2",
  2317 => x"b7c7487e",
  2318 => x"cbc003a8",
  2319 => x"c1486e87",
  2320 => x"c5f1c280",
  2321 => x"87c2c058",
  2322 => x"4dc14cfe",
  2323 => x"ff49fdc3",
  2324 => x"7087f9db",
  2325 => x"0299c249",
  2326 => x"f1c287d5",
  2327 => x"c002bfc1",
  2328 => x"f1c287c9",
  2329 => x"78c048c1",
  2330 => x"fd87c2c0",
  2331 => x"c34dc14c",
  2332 => x"dbff49fa",
  2333 => x"497087d6",
  2334 => x"c00299c2",
  2335 => x"f1c287d9",
  2336 => x"c748bfc1",
  2337 => x"c003a8b7",
  2338 => x"f1c287c9",
  2339 => x"78c748c1",
  2340 => x"fc87c2c0",
  2341 => x"c04dc14c",
  2342 => x"c003acb7",
  2343 => x"66c487d1",
  2344 => x"82d8c14a",
  2345 => x"c6c0026a",
  2346 => x"744b6a87",
  2347 => x"c00f7349",
  2348 => x"1ef0c31e",
  2349 => x"f749dac1",
  2350 => x"86c887d2",
  2351 => x"c0029870",
  2352 => x"a6c887e2",
  2353 => x"c1f1c248",
  2354 => x"66c878bf",
  2355 => x"c491cb49",
  2356 => x"80714866",
  2357 => x"bf6e7e70",
  2358 => x"87c8c002",
  2359 => x"c84bbf6e",
  2360 => x"0f734966",
  2361 => x"c0029d75",
  2362 => x"f1c287c8",
  2363 => x"f349bfc1",
  2364 => x"d5c287c0",
  2365 => x"c002bff5",
  2366 => x"c24987dd",
  2367 => x"987087c7",
  2368 => x"87d3c002",
  2369 => x"bfc1f1c2",
  2370 => x"87e6f249",
  2371 => x"c6f449c0",
  2372 => x"f5d5c287",
  2373 => x"f478c048",
  2374 => x"87e0f38e",
  2375 => x"5c5b5e0e",
  2376 => x"711e0e5d",
  2377 => x"fdf0c24c",
  2378 => x"cdc149bf",
  2379 => x"d1c14da1",
  2380 => x"747e6981",
  2381 => x"87cf029c",
  2382 => x"744ba5c4",
  2383 => x"fdf0c27b",
  2384 => x"fff249bf",
  2385 => x"747b6e87",
  2386 => x"87c4059c",
  2387 => x"87c24bc0",
  2388 => x"49734bc1",
  2389 => x"d487c0f3",
  2390 => x"87c70266",
  2391 => x"7087da49",
  2392 => x"c087c24a",
  2393 => x"f9d5c24a",
  2394 => x"cff2265a",
  2395 => x"00000087",
  2396 => x"00000000",
  2397 => x"00000000",
  2398 => x"4a711e00",
  2399 => x"49bfc8ff",
  2400 => x"2648a172",
  2401 => x"c8ff1e4f",
  2402 => x"c0fe89bf",
  2403 => x"c0c0c0c0",
  2404 => x"87c401a9",
  2405 => x"87c24ac0",
  2406 => x"48724ac1",
  2407 => x"5e0e4f26",
  2408 => x"0e5d5c5b",
  2409 => x"d4ff4b71",
  2410 => x"4866d04c",
  2411 => x"49d678c0",
  2412 => x"87d0d8ff",
  2413 => x"6c7cffc3",
  2414 => x"99ffc349",
  2415 => x"c3494d71",
  2416 => x"e0c199f0",
  2417 => x"87cb05a9",
  2418 => x"6c7cffc3",
  2419 => x"d098c348",
  2420 => x"c3780866",
  2421 => x"4a6c7cff",
  2422 => x"c331c849",
  2423 => x"4a6c7cff",
  2424 => x"4972b271",
  2425 => x"ffc331c8",
  2426 => x"714a6c7c",
  2427 => x"c84972b2",
  2428 => x"7cffc331",
  2429 => x"b2714a6c",
  2430 => x"c048d0ff",
  2431 => x"9b7378e0",
  2432 => x"7287c202",
  2433 => x"2648757b",
  2434 => x"264c264d",
  2435 => x"1e4f264b",
  2436 => x"5e0e4f26",
  2437 => x"f80e5c5b",
  2438 => x"c81e7686",
  2439 => x"fdfd49a6",
  2440 => x"7086c487",
  2441 => x"c2486e4b",
  2442 => x"f0c203a8",
  2443 => x"c34a7387",
  2444 => x"d0c19af0",
  2445 => x"87c702aa",
  2446 => x"05aae0c1",
  2447 => x"7387dec2",
  2448 => x"0299c849",
  2449 => x"c6ff87c3",
  2450 => x"c34c7387",
  2451 => x"05acc29c",
  2452 => x"c487c2c1",
  2453 => x"31c94966",
  2454 => x"66c41e71",
  2455 => x"c292d44a",
  2456 => x"7249c5f1",
  2457 => x"f7cdfe81",
  2458 => x"ff49d887",
  2459 => x"c887d5d5",
  2460 => x"dfc21ec0",
  2461 => x"e9fd49de",
  2462 => x"d0ff87f2",
  2463 => x"78e0c048",
  2464 => x"1ededfc2",
  2465 => x"d44a66cc",
  2466 => x"c5f1c292",
  2467 => x"fe817249",
  2468 => x"cc87fecb",
  2469 => x"05acc186",
  2470 => x"c487c2c1",
  2471 => x"31c94966",
  2472 => x"66c41e71",
  2473 => x"c292d44a",
  2474 => x"7249c5f1",
  2475 => x"efccfe81",
  2476 => x"dedfc287",
  2477 => x"4a66c81e",
  2478 => x"f1c292d4",
  2479 => x"817249c5",
  2480 => x"87fec9fe",
  2481 => x"d3ff49d7",
  2482 => x"c0c887fa",
  2483 => x"dedfc21e",
  2484 => x"f0e7fd49",
  2485 => x"ff86cc87",
  2486 => x"e0c048d0",
  2487 => x"fc8ef878",
  2488 => x"5e0e87e7",
  2489 => x"0e5d5c5b",
  2490 => x"ff4d711e",
  2491 => x"66d44cd4",
  2492 => x"b7c3487e",
  2493 => x"87c506a8",
  2494 => x"e2c148c0",
  2495 => x"fe497587",
  2496 => x"7587c3db",
  2497 => x"4b66c41e",
  2498 => x"f1c293d4",
  2499 => x"497383c5",
  2500 => x"87fac3fe",
  2501 => x"4b6b83c8",
  2502 => x"c848d0ff",
  2503 => x"7cdd78e1",
  2504 => x"ffc34973",
  2505 => x"737c7199",
  2506 => x"29b7c849",
  2507 => x"7199ffc3",
  2508 => x"d049737c",
  2509 => x"ffc329b7",
  2510 => x"737c7199",
  2511 => x"29b7d849",
  2512 => x"7cc07c71",
  2513 => x"7c7c7c7c",
  2514 => x"7c7c7c7c",
  2515 => x"c07c7c7c",
  2516 => x"66c478e0",
  2517 => x"ff49dc1e",
  2518 => x"c887ced2",
  2519 => x"26487386",
  2520 => x"1e87e4fa",
  2521 => x"bff1dec2",
  2522 => x"c2b9c149",
  2523 => x"ff59f5de",
  2524 => x"ffc348d4",
  2525 => x"48d0ff78",
  2526 => x"ff78e1c0",
  2527 => x"78c148d4",
  2528 => x"787131c4",
  2529 => x"c048d0ff",
  2530 => x"4f2678e0",
  2531 => x"e5dec21e",
  2532 => x"d4ecc21e",
  2533 => x"f5c1fe49",
  2534 => x"7086c487",
  2535 => x"87c30298",
  2536 => x"2687c0ff",
  2537 => x"4b35314f",
  2538 => x"20205a48",
  2539 => x"47464320",
  2540 => x"00000000",
  2541 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
