
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"7f",x"00",x"00",x"40"),
     1 => (x"7f",x"19",x"09",x"7f"),
     2 => (x"26",x"00",x"00",x"66"),
     3 => (x"7b",x"59",x"4d",x"6f"),
     4 => (x"01",x"00",x"00",x"32"),
     5 => (x"01",x"7f",x"7f",x"01"),
     6 => (x"3f",x"00",x"00",x"01"),
     7 => (x"7f",x"40",x"40",x"7f"),
     8 => (x"0f",x"00",x"00",x"3f"),
     9 => (x"3f",x"70",x"70",x"3f"),
    10 => (x"7f",x"7f",x"00",x"0f"),
    11 => (x"7f",x"30",x"18",x"30"),
    12 => (x"63",x"41",x"00",x"7f"),
    13 => (x"36",x"1c",x"1c",x"36"),
    14 => (x"03",x"01",x"41",x"63"),
    15 => (x"06",x"7c",x"7c",x"06"),
    16 => (x"71",x"61",x"01",x"03"),
    17 => (x"43",x"47",x"4d",x"59"),
    18 => (x"00",x"00",x"00",x"41"),
    19 => (x"41",x"41",x"7f",x"7f"),
    20 => (x"03",x"01",x"00",x"00"),
    21 => (x"30",x"18",x"0c",x"06"),
    22 => (x"00",x"00",x"40",x"60"),
    23 => (x"7f",x"7f",x"41",x"41"),
    24 => (x"0c",x"08",x"00",x"00"),
    25 => (x"0c",x"06",x"03",x"06"),
    26 => (x"80",x"80",x"00",x"08"),
    27 => (x"80",x"80",x"80",x"80"),
    28 => (x"00",x"00",x"00",x"80"),
    29 => (x"04",x"07",x"03",x"00"),
    30 => (x"20",x"00",x"00",x"00"),
    31 => (x"7c",x"54",x"54",x"74"),
    32 => (x"7f",x"00",x"00",x"78"),
    33 => (x"7c",x"44",x"44",x"7f"),
    34 => (x"38",x"00",x"00",x"38"),
    35 => (x"44",x"44",x"44",x"7c"),
    36 => (x"38",x"00",x"00",x"00"),
    37 => (x"7f",x"44",x"44",x"7c"),
    38 => (x"38",x"00",x"00",x"7f"),
    39 => (x"5c",x"54",x"54",x"7c"),
    40 => (x"04",x"00",x"00",x"18"),
    41 => (x"05",x"05",x"7f",x"7e"),
    42 => (x"18",x"00",x"00",x"00"),
    43 => (x"fc",x"a4",x"a4",x"bc"),
    44 => (x"7f",x"00",x"00",x"7c"),
    45 => (x"7c",x"04",x"04",x"7f"),
    46 => (x"00",x"00",x"00",x"78"),
    47 => (x"40",x"7d",x"3d",x"00"),
    48 => (x"80",x"00",x"00",x"00"),
    49 => (x"7d",x"fd",x"80",x"80"),
    50 => (x"7f",x"00",x"00",x"00"),
    51 => (x"6c",x"38",x"10",x"7f"),
    52 => (x"00",x"00",x"00",x"44"),
    53 => (x"40",x"7f",x"3f",x"00"),
    54 => (x"7c",x"7c",x"00",x"00"),
    55 => (x"7c",x"0c",x"18",x"0c"),
    56 => (x"7c",x"00",x"00",x"78"),
    57 => (x"7c",x"04",x"04",x"7c"),
    58 => (x"38",x"00",x"00",x"78"),
    59 => (x"7c",x"44",x"44",x"7c"),
    60 => (x"fc",x"00",x"00",x"38"),
    61 => (x"3c",x"24",x"24",x"fc"),
    62 => (x"18",x"00",x"00",x"18"),
    63 => (x"fc",x"24",x"24",x"3c"),
    64 => (x"7c",x"00",x"00",x"fc"),
    65 => (x"0c",x"04",x"04",x"7c"),
    66 => (x"48",x"00",x"00",x"08"),
    67 => (x"74",x"54",x"54",x"5c"),
    68 => (x"04",x"00",x"00",x"20"),
    69 => (x"44",x"44",x"7f",x"3f"),
    70 => (x"3c",x"00",x"00",x"00"),
    71 => (x"7c",x"40",x"40",x"7c"),
    72 => (x"1c",x"00",x"00",x"7c"),
    73 => (x"3c",x"60",x"60",x"3c"),
    74 => (x"7c",x"3c",x"00",x"1c"),
    75 => (x"7c",x"60",x"30",x"60"),
    76 => (x"6c",x"44",x"00",x"3c"),
    77 => (x"6c",x"38",x"10",x"38"),
    78 => (x"1c",x"00",x"00",x"44"),
    79 => (x"3c",x"60",x"e0",x"bc"),
    80 => (x"44",x"00",x"00",x"1c"),
    81 => (x"4c",x"5c",x"74",x"64"),
    82 => (x"08",x"00",x"00",x"44"),
    83 => (x"41",x"77",x"3e",x"08"),
    84 => (x"00",x"00",x"00",x"41"),
    85 => (x"00",x"7f",x"7f",x"00"),
    86 => (x"41",x"00",x"00",x"00"),
    87 => (x"08",x"3e",x"77",x"41"),
    88 => (x"01",x"02",x"00",x"08"),
    89 => (x"02",x"02",x"03",x"01"),
    90 => (x"7f",x"7f",x"00",x"01"),
    91 => (x"7f",x"7f",x"7f",x"7f"),
    92 => (x"08",x"08",x"00",x"7f"),
    93 => (x"3e",x"3e",x"1c",x"1c"),
    94 => (x"7f",x"7f",x"7f",x"7f"),
    95 => (x"1c",x"1c",x"3e",x"3e"),
    96 => (x"10",x"00",x"08",x"08"),
    97 => (x"18",x"7c",x"7c",x"18"),
    98 => (x"10",x"00",x"00",x"10"),
    99 => (x"30",x"7c",x"7c",x"30"),
   100 => (x"30",x"10",x"00",x"10"),
   101 => (x"1e",x"78",x"60",x"60"),
   102 => (x"66",x"42",x"00",x"06"),
   103 => (x"66",x"3c",x"18",x"3c"),
   104 => (x"38",x"78",x"00",x"42"),
   105 => (x"6c",x"c6",x"c2",x"6a"),
   106 => (x"00",x"60",x"00",x"38"),
   107 => (x"00",x"00",x"60",x"00"),
   108 => (x"5e",x"0e",x"00",x"60"),
   109 => (x"0e",x"5d",x"5c",x"5b"),
   110 => (x"c2",x"4c",x"71",x"1e"),
   111 => (x"4d",x"bf",x"fd",x"f0"),
   112 => (x"1e",x"c0",x"4b",x"c0"),
   113 => (x"c7",x"02",x"ab",x"74"),
   114 => (x"48",x"a6",x"c4",x"87"),
   115 => (x"87",x"c5",x"78",x"c0"),
   116 => (x"c1",x"48",x"a6",x"c4"),
   117 => (x"1e",x"66",x"c4",x"78"),
   118 => (x"df",x"ee",x"49",x"73"),
   119 => (x"c0",x"86",x"c8",x"87"),
   120 => (x"ef",x"ef",x"49",x"e0"),
   121 => (x"4a",x"a5",x"c4",x"87"),
   122 => (x"f0",x"f0",x"49",x"6a"),
   123 => (x"87",x"c6",x"f1",x"87"),
   124 => (x"83",x"c1",x"85",x"cb"),
   125 => (x"04",x"ab",x"b7",x"c8"),
   126 => (x"26",x"87",x"c7",x"ff"),
   127 => (x"4c",x"26",x"4d",x"26"),
   128 => (x"4f",x"26",x"4b",x"26"),
   129 => (x"c2",x"4a",x"71",x"1e"),
   130 => (x"c2",x"5a",x"c1",x"f1"),
   131 => (x"c7",x"48",x"c1",x"f1"),
   132 => (x"dd",x"fe",x"49",x"78"),
   133 => (x"1e",x"4f",x"26",x"87"),
   134 => (x"4a",x"71",x"1e",x"73"),
   135 => (x"03",x"aa",x"b7",x"c0"),
   136 => (x"d5",x"c2",x"87",x"d3"),
   137 => (x"c4",x"05",x"bf",x"f1"),
   138 => (x"c2",x"4b",x"c1",x"87"),
   139 => (x"c2",x"4b",x"c0",x"87"),
   140 => (x"c4",x"5b",x"f5",x"d5"),
   141 => (x"f5",x"d5",x"c2",x"87"),
   142 => (x"f1",x"d5",x"c2",x"5a"),
   143 => (x"9a",x"c1",x"4a",x"bf"),
   144 => (x"49",x"a2",x"c0",x"c1"),
   145 => (x"fc",x"87",x"e8",x"ec"),
   146 => (x"f1",x"d5",x"c2",x"48"),
   147 => (x"ef",x"fe",x"78",x"bf"),
   148 => (x"4a",x"71",x"1e",x"87"),
   149 => (x"72",x"1e",x"66",x"c4"),
   150 => (x"87",x"e2",x"e6",x"49"),
   151 => (x"1e",x"4f",x"26",x"26"),
   152 => (x"bf",x"f1",x"d5",x"c2"),
   153 => (x"87",x"c4",x"e3",x"49"),
   154 => (x"48",x"f5",x"f0",x"c2"),
   155 => (x"c2",x"78",x"bf",x"e8"),
   156 => (x"ec",x"48",x"f1",x"f0"),
   157 => (x"f0",x"c2",x"78",x"bf"),
   158 => (x"49",x"4a",x"bf",x"f5"),
   159 => (x"c8",x"99",x"ff",x"c3"),
   160 => (x"48",x"72",x"2a",x"b7"),
   161 => (x"f0",x"c2",x"b0",x"71"),
   162 => (x"4f",x"26",x"58",x"fd"),
   163 => (x"5c",x"5b",x"5e",x"0e"),
   164 => (x"4b",x"71",x"0e",x"5d"),
   165 => (x"c2",x"87",x"c8",x"ff"),
   166 => (x"c0",x"48",x"f0",x"f0"),
   167 => (x"e2",x"49",x"73",x"50"),
   168 => (x"49",x"70",x"87",x"ea"),
   169 => (x"cb",x"9c",x"c2",x"4c"),
   170 => (x"cc",x"cb",x"49",x"ee"),
   171 => (x"4d",x"49",x"70",x"87"),
   172 => (x"97",x"f0",x"f0",x"c2"),
   173 => (x"e2",x"c1",x"05",x"bf"),
   174 => (x"49",x"66",x"d0",x"87"),
   175 => (x"bf",x"f9",x"f0",x"c2"),
   176 => (x"87",x"d6",x"05",x"99"),
   177 => (x"c2",x"49",x"66",x"d4"),
   178 => (x"99",x"bf",x"f1",x"f0"),
   179 => (x"73",x"87",x"cb",x"05"),
   180 => (x"87",x"f8",x"e1",x"49"),
   181 => (x"c1",x"02",x"98",x"70"),
   182 => (x"4c",x"c1",x"87",x"c1"),
   183 => (x"75",x"87",x"c0",x"fe"),
   184 => (x"87",x"e1",x"ca",x"49"),
   185 => (x"c6",x"02",x"98",x"70"),
   186 => (x"f0",x"f0",x"c2",x"87"),
   187 => (x"c2",x"50",x"c1",x"48"),
   188 => (x"bf",x"97",x"f0",x"f0"),
   189 => (x"87",x"e3",x"c0",x"05"),
   190 => (x"bf",x"f9",x"f0",x"c2"),
   191 => (x"99",x"66",x"d0",x"49"),
   192 => (x"87",x"d6",x"ff",x"05"),
   193 => (x"bf",x"f1",x"f0",x"c2"),
   194 => (x"99",x"66",x"d4",x"49"),
   195 => (x"87",x"ca",x"ff",x"05"),
   196 => (x"f7",x"e0",x"49",x"73"),
   197 => (x"05",x"98",x"70",x"87"),
   198 => (x"74",x"87",x"ff",x"fe"),
   199 => (x"87",x"dc",x"fb",x"48"),
   200 => (x"5c",x"5b",x"5e",x"0e"),
   201 => (x"86",x"f4",x"0e",x"5d"),
   202 => (x"ec",x"4c",x"4d",x"c0"),
   203 => (x"a6",x"c4",x"7e",x"bf"),
   204 => (x"fd",x"f0",x"c2",x"48"),
   205 => (x"1e",x"c1",x"78",x"bf"),
   206 => (x"49",x"c7",x"1e",x"c0"),
   207 => (x"c8",x"87",x"cd",x"fd"),
   208 => (x"02",x"98",x"70",x"86"),
   209 => (x"49",x"ff",x"87",x"ce"),
   210 => (x"c1",x"87",x"cc",x"fb"),
   211 => (x"df",x"ff",x"49",x"da"),
   212 => (x"4d",x"c1",x"87",x"fa"),
   213 => (x"97",x"f0",x"f0",x"c2"),
   214 => (x"87",x"c3",x"02",x"bf"),
   215 => (x"c2",x"87",x"c4",x"d0"),
   216 => (x"4b",x"bf",x"f5",x"f0"),
   217 => (x"bf",x"f1",x"d5",x"c2"),
   218 => (x"87",x"eb",x"c0",x"05"),
   219 => (x"ff",x"49",x"fd",x"c3"),
   220 => (x"c3",x"87",x"d9",x"df"),
   221 => (x"df",x"ff",x"49",x"fa"),
   222 => (x"49",x"73",x"87",x"d2"),
   223 => (x"71",x"99",x"ff",x"c3"),
   224 => (x"fb",x"49",x"c0",x"1e"),
   225 => (x"49",x"73",x"87",x"cb"),
   226 => (x"71",x"29",x"b7",x"c8"),
   227 => (x"fa",x"49",x"c1",x"1e"),
   228 => (x"86",x"c8",x"87",x"ff"),
   229 => (x"c2",x"87",x"c0",x"c6"),
   230 => (x"4b",x"bf",x"f9",x"f0"),
   231 => (x"87",x"dd",x"02",x"9b"),
   232 => (x"bf",x"ed",x"d5",x"c2"),
   233 => (x"87",x"dd",x"c7",x"49"),
   234 => (x"c4",x"05",x"98",x"70"),
   235 => (x"d2",x"4b",x"c0",x"87"),
   236 => (x"49",x"e0",x"c2",x"87"),
   237 => (x"c2",x"87",x"c2",x"c7"),
   238 => (x"c6",x"58",x"f1",x"d5"),
   239 => (x"ed",x"d5",x"c2",x"87"),
   240 => (x"73",x"78",x"c0",x"48"),
   241 => (x"05",x"99",x"c2",x"49"),
   242 => (x"eb",x"c3",x"87",x"ce"),
   243 => (x"fb",x"dd",x"ff",x"49"),
   244 => (x"c2",x"49",x"70",x"87"),
   245 => (x"87",x"c2",x"02",x"99"),
   246 => (x"49",x"73",x"4c",x"fb"),
   247 => (x"ce",x"05",x"99",x"c1"),
   248 => (x"49",x"f4",x"c3",x"87"),
   249 => (x"87",x"e4",x"dd",x"ff"),
   250 => (x"99",x"c2",x"49",x"70"),
   251 => (x"fa",x"87",x"c2",x"02"),
   252 => (x"c8",x"49",x"73",x"4c"),
   253 => (x"87",x"ce",x"05",x"99"),
   254 => (x"ff",x"49",x"f5",x"c3"),
   255 => (x"70",x"87",x"cd",x"dd"),
   256 => (x"02",x"99",x"c2",x"49"),
   257 => (x"f1",x"c2",x"87",x"d5"),
   258 => (x"ca",x"02",x"bf",x"c1"),
   259 => (x"88",x"c1",x"48",x"87"),
   260 => (x"58",x"c5",x"f1",x"c2"),
   261 => (x"ff",x"87",x"c2",x"c0"),
   262 => (x"73",x"4d",x"c1",x"4c"),
   263 => (x"05",x"99",x"c4",x"49"),
   264 => (x"f2",x"c3",x"87",x"ce"),
   265 => (x"e3",x"dc",x"ff",x"49"),
   266 => (x"c2",x"49",x"70",x"87"),
   267 => (x"87",x"dc",x"02",x"99"),
   268 => (x"bf",x"c1",x"f1",x"c2"),
   269 => (x"b7",x"c7",x"48",x"7e"),
   270 => (x"cb",x"c0",x"03",x"a8"),
   271 => (x"c1",x"48",x"6e",x"87"),
   272 => (x"c5",x"f1",x"c2",x"80"),
   273 => (x"87",x"c2",x"c0",x"58"),
   274 => (x"4d",x"c1",x"4c",x"fe"),
   275 => (x"ff",x"49",x"fd",x"c3"),
   276 => (x"70",x"87",x"f9",x"db"),
   277 => (x"02",x"99",x"c2",x"49"),
   278 => (x"f1",x"c2",x"87",x"d5"),
   279 => (x"c0",x"02",x"bf",x"c1"),
   280 => (x"f1",x"c2",x"87",x"c9"),
   281 => (x"78",x"c0",x"48",x"c1"),
   282 => (x"fd",x"87",x"c2",x"c0"),
   283 => (x"c3",x"4d",x"c1",x"4c"),
   284 => (x"db",x"ff",x"49",x"fa"),
   285 => (x"49",x"70",x"87",x"d6"),
   286 => (x"c0",x"02",x"99",x"c2"),
   287 => (x"f1",x"c2",x"87",x"d9"),
   288 => (x"c7",x"48",x"bf",x"c1"),
   289 => (x"c0",x"03",x"a8",x"b7"),
   290 => (x"f1",x"c2",x"87",x"c9"),
   291 => (x"78",x"c7",x"48",x"c1"),
   292 => (x"fc",x"87",x"c2",x"c0"),
   293 => (x"c0",x"4d",x"c1",x"4c"),
   294 => (x"c0",x"03",x"ac",x"b7"),
   295 => (x"66",x"c4",x"87",x"d1"),
   296 => (x"82",x"d8",x"c1",x"4a"),
   297 => (x"c6",x"c0",x"02",x"6a"),
   298 => (x"74",x"4b",x"6a",x"87"),
   299 => (x"c0",x"0f",x"73",x"49"),
   300 => (x"1e",x"f0",x"c3",x"1e"),
   301 => (x"f7",x"49",x"da",x"c1"),
   302 => (x"86",x"c8",x"87",x"d2"),
   303 => (x"c0",x"02",x"98",x"70"),
   304 => (x"a6",x"c8",x"87",x"e2"),
   305 => (x"c1",x"f1",x"c2",x"48"),
   306 => (x"66",x"c8",x"78",x"bf"),
   307 => (x"c4",x"91",x"cb",x"49"),
   308 => (x"80",x"71",x"48",x"66"),
   309 => (x"bf",x"6e",x"7e",x"70"),
   310 => (x"87",x"c8",x"c0",x"02"),
   311 => (x"c8",x"4b",x"bf",x"6e"),
   312 => (x"0f",x"73",x"49",x"66"),
   313 => (x"c0",x"02",x"9d",x"75"),
   314 => (x"f1",x"c2",x"87",x"c8"),
   315 => (x"f3",x"49",x"bf",x"c1"),
   316 => (x"d5",x"c2",x"87",x"c0"),
   317 => (x"c0",x"02",x"bf",x"f5"),
   318 => (x"c2",x"49",x"87",x"dd"),
   319 => (x"98",x"70",x"87",x"c7"),
   320 => (x"87",x"d3",x"c0",x"02"),
   321 => (x"bf",x"c1",x"f1",x"c2"),
   322 => (x"87",x"e6",x"f2",x"49"),
   323 => (x"c6",x"f4",x"49",x"c0"),
   324 => (x"f5",x"d5",x"c2",x"87"),
   325 => (x"f4",x"78",x"c0",x"48"),
   326 => (x"87",x"e0",x"f3",x"8e"),
   327 => (x"5c",x"5b",x"5e",x"0e"),
   328 => (x"71",x"1e",x"0e",x"5d"),
   329 => (x"fd",x"f0",x"c2",x"4c"),
   330 => (x"cd",x"c1",x"49",x"bf"),
   331 => (x"d1",x"c1",x"4d",x"a1"),
   332 => (x"74",x"7e",x"69",x"81"),
   333 => (x"87",x"cf",x"02",x"9c"),
   334 => (x"74",x"4b",x"a5",x"c4"),
   335 => (x"fd",x"f0",x"c2",x"7b"),
   336 => (x"ff",x"f2",x"49",x"bf"),
   337 => (x"74",x"7b",x"6e",x"87"),
   338 => (x"87",x"c4",x"05",x"9c"),
   339 => (x"87",x"c2",x"4b",x"c0"),
   340 => (x"49",x"73",x"4b",x"c1"),
   341 => (x"d4",x"87",x"c0",x"f3"),
   342 => (x"87",x"c7",x"02",x"66"),
   343 => (x"70",x"87",x"da",x"49"),
   344 => (x"c0",x"87",x"c2",x"4a"),
   345 => (x"f9",x"d5",x"c2",x"4a"),
   346 => (x"cf",x"f2",x"26",x"5a"),
   347 => (x"00",x"00",x"00",x"87"),
   348 => (x"00",x"00",x"00",x"00"),
   349 => (x"00",x"00",x"00",x"00"),
   350 => (x"4a",x"71",x"1e",x"00"),
   351 => (x"49",x"bf",x"c8",x"ff"),
   352 => (x"26",x"48",x"a1",x"72"),
   353 => (x"c8",x"ff",x"1e",x"4f"),
   354 => (x"c0",x"fe",x"89",x"bf"),
   355 => (x"c0",x"c0",x"c0",x"c0"),
   356 => (x"87",x"c4",x"01",x"a9"),
   357 => (x"87",x"c2",x"4a",x"c0"),
   358 => (x"48",x"72",x"4a",x"c1"),
   359 => (x"5e",x"0e",x"4f",x"26"),
   360 => (x"0e",x"5d",x"5c",x"5b"),
   361 => (x"d4",x"ff",x"4b",x"71"),
   362 => (x"48",x"66",x"d0",x"4c"),
   363 => (x"49",x"d6",x"78",x"c0"),
   364 => (x"87",x"d0",x"d8",x"ff"),
   365 => (x"6c",x"7c",x"ff",x"c3"),
   366 => (x"99",x"ff",x"c3",x"49"),
   367 => (x"c3",x"49",x"4d",x"71"),
   368 => (x"e0",x"c1",x"99",x"f0"),
   369 => (x"87",x"cb",x"05",x"a9"),
   370 => (x"6c",x"7c",x"ff",x"c3"),
   371 => (x"d0",x"98",x"c3",x"48"),
   372 => (x"c3",x"78",x"08",x"66"),
   373 => (x"4a",x"6c",x"7c",x"ff"),
   374 => (x"c3",x"31",x"c8",x"49"),
   375 => (x"4a",x"6c",x"7c",x"ff"),
   376 => (x"49",x"72",x"b2",x"71"),
   377 => (x"ff",x"c3",x"31",x"c8"),
   378 => (x"71",x"4a",x"6c",x"7c"),
   379 => (x"c8",x"49",x"72",x"b2"),
   380 => (x"7c",x"ff",x"c3",x"31"),
   381 => (x"b2",x"71",x"4a",x"6c"),
   382 => (x"c0",x"48",x"d0",x"ff"),
   383 => (x"9b",x"73",x"78",x"e0"),
   384 => (x"72",x"87",x"c2",x"02"),
   385 => (x"26",x"48",x"75",x"7b"),
   386 => (x"26",x"4c",x"26",x"4d"),
   387 => (x"1e",x"4f",x"26",x"4b"),
   388 => (x"5e",x"0e",x"4f",x"26"),
   389 => (x"f8",x"0e",x"5c",x"5b"),
   390 => (x"c8",x"1e",x"76",x"86"),
   391 => (x"fd",x"fd",x"49",x"a6"),
   392 => (x"70",x"86",x"c4",x"87"),
   393 => (x"c2",x"48",x"6e",x"4b"),
   394 => (x"f0",x"c2",x"03",x"a8"),
   395 => (x"c3",x"4a",x"73",x"87"),
   396 => (x"d0",x"c1",x"9a",x"f0"),
   397 => (x"87",x"c7",x"02",x"aa"),
   398 => (x"05",x"aa",x"e0",x"c1"),
   399 => (x"73",x"87",x"de",x"c2"),
   400 => (x"02",x"99",x"c8",x"49"),
   401 => (x"c6",x"ff",x"87",x"c3"),
   402 => (x"c3",x"4c",x"73",x"87"),
   403 => (x"05",x"ac",x"c2",x"9c"),
   404 => (x"c4",x"87",x"c2",x"c1"),
   405 => (x"31",x"c9",x"49",x"66"),
   406 => (x"66",x"c4",x"1e",x"71"),
   407 => (x"c2",x"92",x"d4",x"4a"),
   408 => (x"72",x"49",x"c5",x"f1"),
   409 => (x"f7",x"cd",x"fe",x"81"),
   410 => (x"ff",x"49",x"d8",x"87"),
   411 => (x"c8",x"87",x"d5",x"d5"),
   412 => (x"df",x"c2",x"1e",x"c0"),
   413 => (x"e9",x"fd",x"49",x"de"),
   414 => (x"d0",x"ff",x"87",x"f2"),
   415 => (x"78",x"e0",x"c0",x"48"),
   416 => (x"1e",x"de",x"df",x"c2"),
   417 => (x"d4",x"4a",x"66",x"cc"),
   418 => (x"c5",x"f1",x"c2",x"92"),
   419 => (x"fe",x"81",x"72",x"49"),
   420 => (x"cc",x"87",x"fe",x"cb"),
   421 => (x"05",x"ac",x"c1",x"86"),
   422 => (x"c4",x"87",x"c2",x"c1"),
   423 => (x"31",x"c9",x"49",x"66"),
   424 => (x"66",x"c4",x"1e",x"71"),
   425 => (x"c2",x"92",x"d4",x"4a"),
   426 => (x"72",x"49",x"c5",x"f1"),
   427 => (x"ef",x"cc",x"fe",x"81"),
   428 => (x"de",x"df",x"c2",x"87"),
   429 => (x"4a",x"66",x"c8",x"1e"),
   430 => (x"f1",x"c2",x"92",x"d4"),
   431 => (x"81",x"72",x"49",x"c5"),
   432 => (x"87",x"fe",x"c9",x"fe"),
   433 => (x"d3",x"ff",x"49",x"d7"),
   434 => (x"c0",x"c8",x"87",x"fa"),
   435 => (x"de",x"df",x"c2",x"1e"),
   436 => (x"f0",x"e7",x"fd",x"49"),
   437 => (x"ff",x"86",x"cc",x"87"),
   438 => (x"e0",x"c0",x"48",x"d0"),
   439 => (x"fc",x"8e",x"f8",x"78"),
   440 => (x"5e",x"0e",x"87",x"e7"),
   441 => (x"0e",x"5d",x"5c",x"5b"),
   442 => (x"ff",x"4d",x"71",x"1e"),
   443 => (x"66",x"d4",x"4c",x"d4"),
   444 => (x"b7",x"c3",x"48",x"7e"),
   445 => (x"87",x"c5",x"06",x"a8"),
   446 => (x"e2",x"c1",x"48",x"c0"),
   447 => (x"fe",x"49",x"75",x"87"),
   448 => (x"75",x"87",x"c3",x"db"),
   449 => (x"4b",x"66",x"c4",x"1e"),
   450 => (x"f1",x"c2",x"93",x"d4"),
   451 => (x"49",x"73",x"83",x"c5"),
   452 => (x"87",x"fa",x"c3",x"fe"),
   453 => (x"4b",x"6b",x"83",x"c8"),
   454 => (x"c8",x"48",x"d0",x"ff"),
   455 => (x"7c",x"dd",x"78",x"e1"),
   456 => (x"ff",x"c3",x"49",x"73"),
   457 => (x"73",x"7c",x"71",x"99"),
   458 => (x"29",x"b7",x"c8",x"49"),
   459 => (x"71",x"99",x"ff",x"c3"),
   460 => (x"d0",x"49",x"73",x"7c"),
   461 => (x"ff",x"c3",x"29",x"b7"),
   462 => (x"73",x"7c",x"71",x"99"),
   463 => (x"29",x"b7",x"d8",x"49"),
   464 => (x"7c",x"c0",x"7c",x"71"),
   465 => (x"7c",x"7c",x"7c",x"7c"),
   466 => (x"7c",x"7c",x"7c",x"7c"),
   467 => (x"c0",x"7c",x"7c",x"7c"),
   468 => (x"66",x"c4",x"78",x"e0"),
   469 => (x"ff",x"49",x"dc",x"1e"),
   470 => (x"c8",x"87",x"ce",x"d2"),
   471 => (x"26",x"48",x"73",x"86"),
   472 => (x"1e",x"87",x"e4",x"fa"),
   473 => (x"bf",x"f1",x"de",x"c2"),
   474 => (x"c2",x"b9",x"c1",x"49"),
   475 => (x"ff",x"59",x"f5",x"de"),
   476 => (x"ff",x"c3",x"48",x"d4"),
   477 => (x"48",x"d0",x"ff",x"78"),
   478 => (x"ff",x"78",x"e1",x"c0"),
   479 => (x"78",x"c1",x"48",x"d4"),
   480 => (x"78",x"71",x"31",x"c4"),
   481 => (x"c0",x"48",x"d0",x"ff"),
   482 => (x"4f",x"26",x"78",x"e0"),
   483 => (x"e5",x"de",x"c2",x"1e"),
   484 => (x"d4",x"ec",x"c2",x"1e"),
   485 => (x"f5",x"c1",x"fe",x"49"),
   486 => (x"70",x"86",x"c4",x"87"),
   487 => (x"87",x"c3",x"02",x"98"),
   488 => (x"26",x"87",x"c0",x"ff"),
   489 => (x"4b",x"35",x"31",x"4f"),
   490 => (x"20",x"20",x"5a",x"48"),
   491 => (x"47",x"46",x"43",x"20"),
   492 => (x"00",x"00",x"00",x"00"),
   493 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

