
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"7f",x"40",x"40",x"60"),
     1 => (x"7f",x"7f",x"00",x"3f"),
     2 => (x"63",x"36",x"1c",x"08"),
     3 => (x"7f",x"00",x"00",x"41"),
     4 => (x"40",x"40",x"40",x"7f"),
     5 => (x"7f",x"7f",x"00",x"40"),
     6 => (x"7f",x"06",x"0c",x"06"),
     7 => (x"7f",x"7f",x"00",x"7f"),
     8 => (x"7f",x"18",x"0c",x"06"),
     9 => (x"3e",x"00",x"00",x"7f"),
    10 => (x"7f",x"41",x"41",x"7f"),
    11 => (x"7f",x"00",x"00",x"3e"),
    12 => (x"0f",x"09",x"09",x"7f"),
    13 => (x"7f",x"3e",x"00",x"06"),
    14 => (x"7e",x"7f",x"61",x"41"),
    15 => (x"7f",x"00",x"00",x"40"),
    16 => (x"7f",x"19",x"09",x"7f"),
    17 => (x"26",x"00",x"00",x"66"),
    18 => (x"7b",x"59",x"4d",x"6f"),
    19 => (x"01",x"00",x"00",x"32"),
    20 => (x"01",x"7f",x"7f",x"01"),
    21 => (x"3f",x"00",x"00",x"01"),
    22 => (x"7f",x"40",x"40",x"7f"),
    23 => (x"0f",x"00",x"00",x"3f"),
    24 => (x"3f",x"70",x"70",x"3f"),
    25 => (x"7f",x"7f",x"00",x"0f"),
    26 => (x"7f",x"30",x"18",x"30"),
    27 => (x"63",x"41",x"00",x"7f"),
    28 => (x"36",x"1c",x"1c",x"36"),
    29 => (x"03",x"01",x"41",x"63"),
    30 => (x"06",x"7c",x"7c",x"06"),
    31 => (x"71",x"61",x"01",x"03"),
    32 => (x"43",x"47",x"4d",x"59"),
    33 => (x"00",x"00",x"00",x"41"),
    34 => (x"41",x"41",x"7f",x"7f"),
    35 => (x"03",x"01",x"00",x"00"),
    36 => (x"30",x"18",x"0c",x"06"),
    37 => (x"00",x"00",x"40",x"60"),
    38 => (x"7f",x"7f",x"41",x"41"),
    39 => (x"0c",x"08",x"00",x"00"),
    40 => (x"0c",x"06",x"03",x"06"),
    41 => (x"80",x"80",x"00",x"08"),
    42 => (x"80",x"80",x"80",x"80"),
    43 => (x"00",x"00",x"00",x"80"),
    44 => (x"04",x"07",x"03",x"00"),
    45 => (x"20",x"00",x"00",x"00"),
    46 => (x"7c",x"54",x"54",x"74"),
    47 => (x"7f",x"00",x"00",x"78"),
    48 => (x"7c",x"44",x"44",x"7f"),
    49 => (x"38",x"00",x"00",x"38"),
    50 => (x"44",x"44",x"44",x"7c"),
    51 => (x"38",x"00",x"00",x"00"),
    52 => (x"7f",x"44",x"44",x"7c"),
    53 => (x"38",x"00",x"00",x"7f"),
    54 => (x"5c",x"54",x"54",x"7c"),
    55 => (x"04",x"00",x"00",x"18"),
    56 => (x"05",x"05",x"7f",x"7e"),
    57 => (x"18",x"00",x"00",x"00"),
    58 => (x"fc",x"a4",x"a4",x"bc"),
    59 => (x"7f",x"00",x"00",x"7c"),
    60 => (x"7c",x"04",x"04",x"7f"),
    61 => (x"00",x"00",x"00",x"78"),
    62 => (x"40",x"7d",x"3d",x"00"),
    63 => (x"80",x"00",x"00",x"00"),
    64 => (x"7d",x"fd",x"80",x"80"),
    65 => (x"7f",x"00",x"00",x"00"),
    66 => (x"6c",x"38",x"10",x"7f"),
    67 => (x"00",x"00",x"00",x"44"),
    68 => (x"40",x"7f",x"3f",x"00"),
    69 => (x"7c",x"7c",x"00",x"00"),
    70 => (x"7c",x"0c",x"18",x"0c"),
    71 => (x"7c",x"00",x"00",x"78"),
    72 => (x"7c",x"04",x"04",x"7c"),
    73 => (x"38",x"00",x"00",x"78"),
    74 => (x"7c",x"44",x"44",x"7c"),
    75 => (x"fc",x"00",x"00",x"38"),
    76 => (x"3c",x"24",x"24",x"fc"),
    77 => (x"18",x"00",x"00",x"18"),
    78 => (x"fc",x"24",x"24",x"3c"),
    79 => (x"7c",x"00",x"00",x"fc"),
    80 => (x"0c",x"04",x"04",x"7c"),
    81 => (x"48",x"00",x"00",x"08"),
    82 => (x"74",x"54",x"54",x"5c"),
    83 => (x"04",x"00",x"00",x"20"),
    84 => (x"44",x"44",x"7f",x"3f"),
    85 => (x"3c",x"00",x"00",x"00"),
    86 => (x"7c",x"40",x"40",x"7c"),
    87 => (x"1c",x"00",x"00",x"7c"),
    88 => (x"3c",x"60",x"60",x"3c"),
    89 => (x"7c",x"3c",x"00",x"1c"),
    90 => (x"7c",x"60",x"30",x"60"),
    91 => (x"6c",x"44",x"00",x"3c"),
    92 => (x"6c",x"38",x"10",x"38"),
    93 => (x"1c",x"00",x"00",x"44"),
    94 => (x"3c",x"60",x"e0",x"bc"),
    95 => (x"44",x"00",x"00",x"1c"),
    96 => (x"4c",x"5c",x"74",x"64"),
    97 => (x"08",x"00",x"00",x"44"),
    98 => (x"41",x"77",x"3e",x"08"),
    99 => (x"00",x"00",x"00",x"41"),
   100 => (x"00",x"7f",x"7f",x"00"),
   101 => (x"41",x"00",x"00",x"00"),
   102 => (x"08",x"3e",x"77",x"41"),
   103 => (x"01",x"02",x"00",x"08"),
   104 => (x"02",x"02",x"03",x"01"),
   105 => (x"7f",x"7f",x"00",x"01"),
   106 => (x"7f",x"7f",x"7f",x"7f"),
   107 => (x"08",x"08",x"00",x"7f"),
   108 => (x"3e",x"3e",x"1c",x"1c"),
   109 => (x"7f",x"7f",x"7f",x"7f"),
   110 => (x"1c",x"1c",x"3e",x"3e"),
   111 => (x"10",x"00",x"08",x"08"),
   112 => (x"18",x"7c",x"7c",x"18"),
   113 => (x"10",x"00",x"00",x"10"),
   114 => (x"30",x"7c",x"7c",x"30"),
   115 => (x"30",x"10",x"00",x"10"),
   116 => (x"1e",x"78",x"60",x"60"),
   117 => (x"66",x"42",x"00",x"06"),
   118 => (x"66",x"3c",x"18",x"3c"),
   119 => (x"38",x"78",x"00",x"42"),
   120 => (x"6c",x"c6",x"c2",x"6a"),
   121 => (x"00",x"60",x"00",x"38"),
   122 => (x"00",x"00",x"60",x"00"),
   123 => (x"5e",x"0e",x"00",x"60"),
   124 => (x"0e",x"5d",x"5c",x"5b"),
   125 => (x"c2",x"4c",x"71",x"1e"),
   126 => (x"4d",x"bf",x"d1",x"f1"),
   127 => (x"1e",x"c0",x"4b",x"c0"),
   128 => (x"c7",x"02",x"ab",x"74"),
   129 => (x"48",x"a6",x"c4",x"87"),
   130 => (x"87",x"c5",x"78",x"c0"),
   131 => (x"c1",x"48",x"a6",x"c4"),
   132 => (x"1e",x"66",x"c4",x"78"),
   133 => (x"df",x"ee",x"49",x"73"),
   134 => (x"c0",x"86",x"c8",x"87"),
   135 => (x"ef",x"ef",x"49",x"e0"),
   136 => (x"4a",x"a5",x"c4",x"87"),
   137 => (x"f0",x"f0",x"49",x"6a"),
   138 => (x"87",x"c6",x"f1",x"87"),
   139 => (x"83",x"c1",x"85",x"cb"),
   140 => (x"04",x"ab",x"b7",x"c8"),
   141 => (x"26",x"87",x"c7",x"ff"),
   142 => (x"4c",x"26",x"4d",x"26"),
   143 => (x"4f",x"26",x"4b",x"26"),
   144 => (x"c2",x"4a",x"71",x"1e"),
   145 => (x"c2",x"5a",x"d5",x"f1"),
   146 => (x"c7",x"48",x"d5",x"f1"),
   147 => (x"dd",x"fe",x"49",x"78"),
   148 => (x"1e",x"4f",x"26",x"87"),
   149 => (x"4a",x"71",x"1e",x"73"),
   150 => (x"03",x"aa",x"b7",x"c0"),
   151 => (x"d6",x"c2",x"87",x"d3"),
   152 => (x"c4",x"05",x"bf",x"ed"),
   153 => (x"c2",x"4b",x"c1",x"87"),
   154 => (x"c2",x"4b",x"c0",x"87"),
   155 => (x"c4",x"5b",x"f1",x"d6"),
   156 => (x"f1",x"d6",x"c2",x"87"),
   157 => (x"ed",x"d6",x"c2",x"5a"),
   158 => (x"9a",x"c1",x"4a",x"bf"),
   159 => (x"49",x"a2",x"c0",x"c1"),
   160 => (x"fc",x"87",x"e8",x"ec"),
   161 => (x"ed",x"d6",x"c2",x"48"),
   162 => (x"ef",x"fe",x"78",x"bf"),
   163 => (x"4a",x"71",x"1e",x"87"),
   164 => (x"72",x"1e",x"66",x"c4"),
   165 => (x"87",x"e2",x"e6",x"49"),
   166 => (x"1e",x"4f",x"26",x"26"),
   167 => (x"bf",x"ed",x"d6",x"c2"),
   168 => (x"87",x"c4",x"e3",x"49"),
   169 => (x"48",x"c9",x"f1",x"c2"),
   170 => (x"c2",x"78",x"bf",x"e8"),
   171 => (x"ec",x"48",x"c5",x"f1"),
   172 => (x"f1",x"c2",x"78",x"bf"),
   173 => (x"49",x"4a",x"bf",x"c9"),
   174 => (x"c8",x"99",x"ff",x"c3"),
   175 => (x"48",x"72",x"2a",x"b7"),
   176 => (x"f1",x"c2",x"b0",x"71"),
   177 => (x"4f",x"26",x"58",x"d1"),
   178 => (x"5c",x"5b",x"5e",x"0e"),
   179 => (x"4b",x"71",x"0e",x"5d"),
   180 => (x"c2",x"87",x"c8",x"ff"),
   181 => (x"c0",x"48",x"c4",x"f1"),
   182 => (x"e2",x"49",x"73",x"50"),
   183 => (x"49",x"70",x"87",x"ea"),
   184 => (x"cb",x"9c",x"c2",x"4c"),
   185 => (x"cc",x"cb",x"49",x"ee"),
   186 => (x"4d",x"49",x"70",x"87"),
   187 => (x"97",x"c4",x"f1",x"c2"),
   188 => (x"e2",x"c1",x"05",x"bf"),
   189 => (x"49",x"66",x"d0",x"87"),
   190 => (x"bf",x"cd",x"f1",x"c2"),
   191 => (x"87",x"d6",x"05",x"99"),
   192 => (x"c2",x"49",x"66",x"d4"),
   193 => (x"99",x"bf",x"c5",x"f1"),
   194 => (x"73",x"87",x"cb",x"05"),
   195 => (x"87",x"f8",x"e1",x"49"),
   196 => (x"c1",x"02",x"98",x"70"),
   197 => (x"4c",x"c1",x"87",x"c1"),
   198 => (x"75",x"87",x"c0",x"fe"),
   199 => (x"87",x"e1",x"ca",x"49"),
   200 => (x"c6",x"02",x"98",x"70"),
   201 => (x"c4",x"f1",x"c2",x"87"),
   202 => (x"c2",x"50",x"c1",x"48"),
   203 => (x"bf",x"97",x"c4",x"f1"),
   204 => (x"87",x"e3",x"c0",x"05"),
   205 => (x"bf",x"cd",x"f1",x"c2"),
   206 => (x"99",x"66",x"d0",x"49"),
   207 => (x"87",x"d6",x"ff",x"05"),
   208 => (x"bf",x"c5",x"f1",x"c2"),
   209 => (x"99",x"66",x"d4",x"49"),
   210 => (x"87",x"ca",x"ff",x"05"),
   211 => (x"f7",x"e0",x"49",x"73"),
   212 => (x"05",x"98",x"70",x"87"),
   213 => (x"74",x"87",x"ff",x"fe"),
   214 => (x"87",x"dc",x"fb",x"48"),
   215 => (x"5c",x"5b",x"5e",x"0e"),
   216 => (x"86",x"f4",x"0e",x"5d"),
   217 => (x"ec",x"4c",x"4d",x"c0"),
   218 => (x"a6",x"c4",x"7e",x"bf"),
   219 => (x"d1",x"f1",x"c2",x"48"),
   220 => (x"1e",x"c1",x"78",x"bf"),
   221 => (x"49",x"c7",x"1e",x"c0"),
   222 => (x"c8",x"87",x"cd",x"fd"),
   223 => (x"02",x"98",x"70",x"86"),
   224 => (x"49",x"ff",x"87",x"ce"),
   225 => (x"c1",x"87",x"cc",x"fb"),
   226 => (x"df",x"ff",x"49",x"da"),
   227 => (x"4d",x"c1",x"87",x"fa"),
   228 => (x"97",x"c4",x"f1",x"c2"),
   229 => (x"87",x"c3",x"02",x"bf"),
   230 => (x"c2",x"87",x"c4",x"d0"),
   231 => (x"4b",x"bf",x"c9",x"f1"),
   232 => (x"bf",x"ed",x"d6",x"c2"),
   233 => (x"87",x"eb",x"c0",x"05"),
   234 => (x"ff",x"49",x"fd",x"c3"),
   235 => (x"c3",x"87",x"d9",x"df"),
   236 => (x"df",x"ff",x"49",x"fa"),
   237 => (x"49",x"73",x"87",x"d2"),
   238 => (x"71",x"99",x"ff",x"c3"),
   239 => (x"fb",x"49",x"c0",x"1e"),
   240 => (x"49",x"73",x"87",x"cb"),
   241 => (x"71",x"29",x"b7",x"c8"),
   242 => (x"fa",x"49",x"c1",x"1e"),
   243 => (x"86",x"c8",x"87",x"ff"),
   244 => (x"c2",x"87",x"c0",x"c6"),
   245 => (x"4b",x"bf",x"cd",x"f1"),
   246 => (x"87",x"dd",x"02",x"9b"),
   247 => (x"bf",x"e9",x"d6",x"c2"),
   248 => (x"87",x"dd",x"c7",x"49"),
   249 => (x"c4",x"05",x"98",x"70"),
   250 => (x"d2",x"4b",x"c0",x"87"),
   251 => (x"49",x"e0",x"c2",x"87"),
   252 => (x"c2",x"87",x"c2",x"c7"),
   253 => (x"c6",x"58",x"ed",x"d6"),
   254 => (x"e9",x"d6",x"c2",x"87"),
   255 => (x"73",x"78",x"c0",x"48"),
   256 => (x"05",x"99",x"c2",x"49"),
   257 => (x"eb",x"c3",x"87",x"ce"),
   258 => (x"fb",x"dd",x"ff",x"49"),
   259 => (x"c2",x"49",x"70",x"87"),
   260 => (x"87",x"c2",x"02",x"99"),
   261 => (x"49",x"73",x"4c",x"fb"),
   262 => (x"ce",x"05",x"99",x"c1"),
   263 => (x"49",x"f4",x"c3",x"87"),
   264 => (x"87",x"e4",x"dd",x"ff"),
   265 => (x"99",x"c2",x"49",x"70"),
   266 => (x"fa",x"87",x"c2",x"02"),
   267 => (x"c8",x"49",x"73",x"4c"),
   268 => (x"87",x"ce",x"05",x"99"),
   269 => (x"ff",x"49",x"f5",x"c3"),
   270 => (x"70",x"87",x"cd",x"dd"),
   271 => (x"02",x"99",x"c2",x"49"),
   272 => (x"f1",x"c2",x"87",x"d5"),
   273 => (x"ca",x"02",x"bf",x"d5"),
   274 => (x"88",x"c1",x"48",x"87"),
   275 => (x"58",x"d9",x"f1",x"c2"),
   276 => (x"ff",x"87",x"c2",x"c0"),
   277 => (x"73",x"4d",x"c1",x"4c"),
   278 => (x"05",x"99",x"c4",x"49"),
   279 => (x"f2",x"c3",x"87",x"ce"),
   280 => (x"e3",x"dc",x"ff",x"49"),
   281 => (x"c2",x"49",x"70",x"87"),
   282 => (x"87",x"dc",x"02",x"99"),
   283 => (x"bf",x"d5",x"f1",x"c2"),
   284 => (x"b7",x"c7",x"48",x"7e"),
   285 => (x"cb",x"c0",x"03",x"a8"),
   286 => (x"c1",x"48",x"6e",x"87"),
   287 => (x"d9",x"f1",x"c2",x"80"),
   288 => (x"87",x"c2",x"c0",x"58"),
   289 => (x"4d",x"c1",x"4c",x"fe"),
   290 => (x"ff",x"49",x"fd",x"c3"),
   291 => (x"70",x"87",x"f9",x"db"),
   292 => (x"02",x"99",x"c2",x"49"),
   293 => (x"f1",x"c2",x"87",x"d5"),
   294 => (x"c0",x"02",x"bf",x"d5"),
   295 => (x"f1",x"c2",x"87",x"c9"),
   296 => (x"78",x"c0",x"48",x"d5"),
   297 => (x"fd",x"87",x"c2",x"c0"),
   298 => (x"c3",x"4d",x"c1",x"4c"),
   299 => (x"db",x"ff",x"49",x"fa"),
   300 => (x"49",x"70",x"87",x"d6"),
   301 => (x"c0",x"02",x"99",x"c2"),
   302 => (x"f1",x"c2",x"87",x"d9"),
   303 => (x"c7",x"48",x"bf",x"d5"),
   304 => (x"c0",x"03",x"a8",x"b7"),
   305 => (x"f1",x"c2",x"87",x"c9"),
   306 => (x"78",x"c7",x"48",x"d5"),
   307 => (x"fc",x"87",x"c2",x"c0"),
   308 => (x"c0",x"4d",x"c1",x"4c"),
   309 => (x"c0",x"03",x"ac",x"b7"),
   310 => (x"66",x"c4",x"87",x"d1"),
   311 => (x"82",x"d8",x"c1",x"4a"),
   312 => (x"c6",x"c0",x"02",x"6a"),
   313 => (x"74",x"4b",x"6a",x"87"),
   314 => (x"c0",x"0f",x"73",x"49"),
   315 => (x"1e",x"f0",x"c3",x"1e"),
   316 => (x"f7",x"49",x"da",x"c1"),
   317 => (x"86",x"c8",x"87",x"d2"),
   318 => (x"c0",x"02",x"98",x"70"),
   319 => (x"a6",x"c8",x"87",x"e2"),
   320 => (x"d5",x"f1",x"c2",x"48"),
   321 => (x"66",x"c8",x"78",x"bf"),
   322 => (x"c4",x"91",x"cb",x"49"),
   323 => (x"80",x"71",x"48",x"66"),
   324 => (x"bf",x"6e",x"7e",x"70"),
   325 => (x"87",x"c8",x"c0",x"02"),
   326 => (x"c8",x"4b",x"bf",x"6e"),
   327 => (x"0f",x"73",x"49",x"66"),
   328 => (x"c0",x"02",x"9d",x"75"),
   329 => (x"f1",x"c2",x"87",x"c8"),
   330 => (x"f3",x"49",x"bf",x"d5"),
   331 => (x"d6",x"c2",x"87",x"c0"),
   332 => (x"c0",x"02",x"bf",x"f1"),
   333 => (x"c2",x"49",x"87",x"dd"),
   334 => (x"98",x"70",x"87",x"c7"),
   335 => (x"87",x"d3",x"c0",x"02"),
   336 => (x"bf",x"d5",x"f1",x"c2"),
   337 => (x"87",x"e6",x"f2",x"49"),
   338 => (x"c6",x"f4",x"49",x"c0"),
   339 => (x"f1",x"d6",x"c2",x"87"),
   340 => (x"f4",x"78",x"c0",x"48"),
   341 => (x"87",x"e0",x"f3",x"8e"),
   342 => (x"5c",x"5b",x"5e",x"0e"),
   343 => (x"71",x"1e",x"0e",x"5d"),
   344 => (x"d1",x"f1",x"c2",x"4c"),
   345 => (x"cd",x"c1",x"49",x"bf"),
   346 => (x"d1",x"c1",x"4d",x"a1"),
   347 => (x"74",x"7e",x"69",x"81"),
   348 => (x"87",x"cf",x"02",x"9c"),
   349 => (x"74",x"4b",x"a5",x"c4"),
   350 => (x"d1",x"f1",x"c2",x"7b"),
   351 => (x"ff",x"f2",x"49",x"bf"),
   352 => (x"74",x"7b",x"6e",x"87"),
   353 => (x"87",x"c4",x"05",x"9c"),
   354 => (x"87",x"c2",x"4b",x"c0"),
   355 => (x"49",x"73",x"4b",x"c1"),
   356 => (x"d4",x"87",x"c0",x"f3"),
   357 => (x"87",x"c7",x"02",x"66"),
   358 => (x"70",x"87",x"da",x"49"),
   359 => (x"c0",x"87",x"c2",x"4a"),
   360 => (x"f5",x"d6",x"c2",x"4a"),
   361 => (x"cf",x"f2",x"26",x"5a"),
   362 => (x"00",x"00",x"00",x"87"),
   363 => (x"00",x"00",x"00",x"00"),
   364 => (x"00",x"00",x"00",x"00"),
   365 => (x"4a",x"71",x"1e",x"00"),
   366 => (x"49",x"bf",x"c8",x"ff"),
   367 => (x"26",x"48",x"a1",x"72"),
   368 => (x"c8",x"ff",x"1e",x"4f"),
   369 => (x"c0",x"fe",x"89",x"bf"),
   370 => (x"c0",x"c0",x"c0",x"c0"),
   371 => (x"87",x"c4",x"01",x"a9"),
   372 => (x"87",x"c2",x"4a",x"c0"),
   373 => (x"48",x"72",x"4a",x"c1"),
   374 => (x"5e",x"0e",x"4f",x"26"),
   375 => (x"0e",x"5d",x"5c",x"5b"),
   376 => (x"d4",x"ff",x"4b",x"71"),
   377 => (x"48",x"66",x"d0",x"4c"),
   378 => (x"49",x"d6",x"78",x"c0"),
   379 => (x"87",x"d0",x"d8",x"ff"),
   380 => (x"6c",x"7c",x"ff",x"c3"),
   381 => (x"99",x"ff",x"c3",x"49"),
   382 => (x"c3",x"49",x"4d",x"71"),
   383 => (x"e0",x"c1",x"99",x"f0"),
   384 => (x"87",x"cb",x"05",x"a9"),
   385 => (x"6c",x"7c",x"ff",x"c3"),
   386 => (x"d0",x"98",x"c3",x"48"),
   387 => (x"c3",x"78",x"08",x"66"),
   388 => (x"4a",x"6c",x"7c",x"ff"),
   389 => (x"c3",x"31",x"c8",x"49"),
   390 => (x"4a",x"6c",x"7c",x"ff"),
   391 => (x"49",x"72",x"b2",x"71"),
   392 => (x"ff",x"c3",x"31",x"c8"),
   393 => (x"71",x"4a",x"6c",x"7c"),
   394 => (x"c8",x"49",x"72",x"b2"),
   395 => (x"7c",x"ff",x"c3",x"31"),
   396 => (x"b2",x"71",x"4a",x"6c"),
   397 => (x"c0",x"48",x"d0",x"ff"),
   398 => (x"9b",x"73",x"78",x"e0"),
   399 => (x"72",x"87",x"c2",x"02"),
   400 => (x"26",x"48",x"75",x"7b"),
   401 => (x"26",x"4c",x"26",x"4d"),
   402 => (x"1e",x"4f",x"26",x"4b"),
   403 => (x"5e",x"0e",x"4f",x"26"),
   404 => (x"f8",x"0e",x"5c",x"5b"),
   405 => (x"c8",x"1e",x"76",x"86"),
   406 => (x"fd",x"fd",x"49",x"a6"),
   407 => (x"70",x"86",x"c4",x"87"),
   408 => (x"c2",x"48",x"6e",x"4b"),
   409 => (x"f0",x"c2",x"03",x"a8"),
   410 => (x"c3",x"4a",x"73",x"87"),
   411 => (x"d0",x"c1",x"9a",x"f0"),
   412 => (x"87",x"c7",x"02",x"aa"),
   413 => (x"05",x"aa",x"e0",x"c1"),
   414 => (x"73",x"87",x"de",x"c2"),
   415 => (x"02",x"99",x"c8",x"49"),
   416 => (x"c6",x"ff",x"87",x"c3"),
   417 => (x"c3",x"4c",x"73",x"87"),
   418 => (x"05",x"ac",x"c2",x"9c"),
   419 => (x"c4",x"87",x"c2",x"c1"),
   420 => (x"31",x"c9",x"49",x"66"),
   421 => (x"66",x"c4",x"1e",x"71"),
   422 => (x"c2",x"92",x"d4",x"4a"),
   423 => (x"72",x"49",x"d9",x"f1"),
   424 => (x"ed",x"cc",x"fe",x"81"),
   425 => (x"ff",x"49",x"d8",x"87"),
   426 => (x"c8",x"87",x"d5",x"d5"),
   427 => (x"df",x"c2",x"1e",x"c0"),
   428 => (x"e8",x"fd",x"49",x"f2"),
   429 => (x"d0",x"ff",x"87",x"e9"),
   430 => (x"78",x"e0",x"c0",x"48"),
   431 => (x"1e",x"f2",x"df",x"c2"),
   432 => (x"d4",x"4a",x"66",x"cc"),
   433 => (x"d9",x"f1",x"c2",x"92"),
   434 => (x"fe",x"81",x"72",x"49"),
   435 => (x"cc",x"87",x"f4",x"ca"),
   436 => (x"05",x"ac",x"c1",x"86"),
   437 => (x"c4",x"87",x"c2",x"c1"),
   438 => (x"31",x"c9",x"49",x"66"),
   439 => (x"66",x"c4",x"1e",x"71"),
   440 => (x"c2",x"92",x"d4",x"4a"),
   441 => (x"72",x"49",x"d9",x"f1"),
   442 => (x"e5",x"cb",x"fe",x"81"),
   443 => (x"f2",x"df",x"c2",x"87"),
   444 => (x"4a",x"66",x"c8",x"1e"),
   445 => (x"f1",x"c2",x"92",x"d4"),
   446 => (x"81",x"72",x"49",x"d9"),
   447 => (x"87",x"f4",x"c8",x"fe"),
   448 => (x"d3",x"ff",x"49",x"d7"),
   449 => (x"c0",x"c8",x"87",x"fa"),
   450 => (x"f2",x"df",x"c2",x"1e"),
   451 => (x"e7",x"e6",x"fd",x"49"),
   452 => (x"ff",x"86",x"cc",x"87"),
   453 => (x"e0",x"c0",x"48",x"d0"),
   454 => (x"fc",x"8e",x"f8",x"78"),
   455 => (x"5e",x"0e",x"87",x"e7"),
   456 => (x"0e",x"5d",x"5c",x"5b"),
   457 => (x"ff",x"4d",x"71",x"1e"),
   458 => (x"66",x"d4",x"4c",x"d4"),
   459 => (x"b7",x"c3",x"48",x"7e"),
   460 => (x"87",x"c5",x"06",x"a8"),
   461 => (x"e2",x"c1",x"48",x"c0"),
   462 => (x"fe",x"49",x"75",x"87"),
   463 => (x"75",x"87",x"f8",x"d9"),
   464 => (x"4b",x"66",x"c4",x"1e"),
   465 => (x"f1",x"c2",x"93",x"d4"),
   466 => (x"49",x"73",x"83",x"d9"),
   467 => (x"87",x"f1",x"c2",x"fe"),
   468 => (x"4b",x"6b",x"83",x"c8"),
   469 => (x"c8",x"48",x"d0",x"ff"),
   470 => (x"7c",x"dd",x"78",x"e1"),
   471 => (x"ff",x"c3",x"49",x"73"),
   472 => (x"73",x"7c",x"71",x"99"),
   473 => (x"29",x"b7",x"c8",x"49"),
   474 => (x"71",x"99",x"ff",x"c3"),
   475 => (x"d0",x"49",x"73",x"7c"),
   476 => (x"ff",x"c3",x"29",x"b7"),
   477 => (x"73",x"7c",x"71",x"99"),
   478 => (x"29",x"b7",x"d8",x"49"),
   479 => (x"7c",x"c0",x"7c",x"71"),
   480 => (x"7c",x"7c",x"7c",x"7c"),
   481 => (x"7c",x"7c",x"7c",x"7c"),
   482 => (x"c0",x"7c",x"7c",x"7c"),
   483 => (x"66",x"c4",x"78",x"e0"),
   484 => (x"ff",x"49",x"dc",x"1e"),
   485 => (x"c8",x"87",x"ce",x"d2"),
   486 => (x"26",x"48",x"73",x"86"),
   487 => (x"1e",x"87",x"e4",x"fa"),
   488 => (x"bf",x"c8",x"df",x"c2"),
   489 => (x"c2",x"b9",x"c1",x"49"),
   490 => (x"ff",x"59",x"cc",x"df"),
   491 => (x"ff",x"c3",x"48",x"d4"),
   492 => (x"48",x"d0",x"ff",x"78"),
   493 => (x"ff",x"78",x"e1",x"c0"),
   494 => (x"78",x"c1",x"48",x"d4"),
   495 => (x"78",x"71",x"31",x"c4"),
   496 => (x"c0",x"48",x"d0",x"ff"),
   497 => (x"4f",x"26",x"78",x"e0"),
   498 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

