package build_id is
constant BUILD_DATE : string := "230424";
constant BUILD_TIME : string := "145844";
end build_id;
