
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f4",x"f1",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"f4",x"f1",x"c2"),
    14 => (x"48",x"fc",x"de",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"dd",x"e1"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"4a",x"71",x"1e",x"4f"),
    50 => (x"48",x"49",x"66",x"c4"),
    51 => (x"a6",x"c8",x"88",x"c1"),
    52 => (x"02",x"99",x"71",x"58"),
    53 => (x"48",x"12",x"87",x"d4"),
    54 => (x"78",x"08",x"d4",x"ff"),
    55 => (x"48",x"49",x"66",x"c4"),
    56 => (x"a6",x"c8",x"88",x"c1"),
    57 => (x"05",x"99",x"71",x"58"),
    58 => (x"4f",x"26",x"87",x"ec"),
    59 => (x"c4",x"4a",x"71",x"1e"),
    60 => (x"c1",x"48",x"49",x"66"),
    61 => (x"58",x"a6",x"c8",x"88"),
    62 => (x"d6",x"02",x"99",x"71"),
    63 => (x"48",x"d4",x"ff",x"87"),
    64 => (x"68",x"78",x"ff",x"c3"),
    65 => (x"49",x"66",x"c4",x"52"),
    66 => (x"c8",x"88",x"c1",x"48"),
    67 => (x"99",x"71",x"58",x"a6"),
    68 => (x"26",x"87",x"ea",x"05"),
    69 => (x"1e",x"73",x"1e",x"4f"),
    70 => (x"c3",x"4b",x"d4",x"ff"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"6b",x"7b",x"ff",x"c3"),
    73 => (x"72",x"32",x"c8",x"49"),
    74 => (x"7b",x"ff",x"c3",x"b1"),
    75 => (x"31",x"c8",x"4a",x"6b"),
    76 => (x"ff",x"c3",x"b2",x"71"),
    77 => (x"c8",x"49",x"6b",x"7b"),
    78 => (x"71",x"b1",x"72",x"32"),
    79 => (x"26",x"87",x"c4",x"48"),
    80 => (x"26",x"4c",x"26",x"4d"),
    81 => (x"0e",x"4f",x"26",x"4b"),
    82 => (x"5d",x"5c",x"5b",x"5e"),
    83 => (x"ff",x"4a",x"71",x"0e"),
    84 => (x"49",x"72",x"4c",x"d4"),
    85 => (x"71",x"99",x"ff",x"c3"),
    86 => (x"fc",x"de",x"c2",x"7c"),
    87 => (x"87",x"c8",x"05",x"bf"),
    88 => (x"c9",x"48",x"66",x"d0"),
    89 => (x"58",x"a6",x"d4",x"30"),
    90 => (x"d8",x"49",x"66",x"d0"),
    91 => (x"99",x"ff",x"c3",x"29"),
    92 => (x"66",x"d0",x"7c",x"71"),
    93 => (x"c3",x"29",x"d0",x"49"),
    94 => (x"7c",x"71",x"99",x"ff"),
    95 => (x"c8",x"49",x"66",x"d0"),
    96 => (x"99",x"ff",x"c3",x"29"),
    97 => (x"66",x"d0",x"7c",x"71"),
    98 => (x"99",x"ff",x"c3",x"49"),
    99 => (x"49",x"72",x"7c",x"71"),
   100 => (x"ff",x"c3",x"29",x"d0"),
   101 => (x"6c",x"7c",x"71",x"99"),
   102 => (x"ff",x"f0",x"c9",x"4b"),
   103 => (x"ab",x"ff",x"c3",x"4d"),
   104 => (x"c3",x"87",x"d0",x"05"),
   105 => (x"4b",x"6c",x"7c",x"ff"),
   106 => (x"c6",x"02",x"8d",x"c1"),
   107 => (x"ab",x"ff",x"c3",x"87"),
   108 => (x"73",x"87",x"f0",x"02"),
   109 => (x"87",x"c7",x"fe",x"48"),
   110 => (x"ff",x"49",x"c0",x"1e"),
   111 => (x"ff",x"c3",x"48",x"d4"),
   112 => (x"c3",x"81",x"c1",x"78"),
   113 => (x"04",x"a9",x"b7",x"c8"),
   114 => (x"4f",x"26",x"87",x"f1"),
   115 => (x"e7",x"1e",x"73",x"1e"),
   116 => (x"df",x"f8",x"c4",x"87"),
   117 => (x"c0",x"1e",x"c0",x"4b"),
   118 => (x"f7",x"c1",x"f0",x"ff"),
   119 => (x"87",x"e7",x"fd",x"49"),
   120 => (x"a8",x"c1",x"86",x"c4"),
   121 => (x"87",x"ea",x"c0",x"05"),
   122 => (x"c3",x"48",x"d4",x"ff"),
   123 => (x"c0",x"c1",x"78",x"ff"),
   124 => (x"c0",x"c0",x"c0",x"c0"),
   125 => (x"f0",x"e1",x"c0",x"1e"),
   126 => (x"fd",x"49",x"e9",x"c1"),
   127 => (x"86",x"c4",x"87",x"c9"),
   128 => (x"ca",x"05",x"98",x"70"),
   129 => (x"48",x"d4",x"ff",x"87"),
   130 => (x"c1",x"78",x"ff",x"c3"),
   131 => (x"fe",x"87",x"cb",x"48"),
   132 => (x"8b",x"c1",x"87",x"e6"),
   133 => (x"87",x"fd",x"fe",x"05"),
   134 => (x"e6",x"fc",x"48",x"c0"),
   135 => (x"1e",x"73",x"1e",x"87"),
   136 => (x"c3",x"48",x"d4",x"ff"),
   137 => (x"4b",x"d3",x"78",x"ff"),
   138 => (x"ff",x"c0",x"1e",x"c0"),
   139 => (x"49",x"c1",x"c1",x"f0"),
   140 => (x"c4",x"87",x"d4",x"fc"),
   141 => (x"05",x"98",x"70",x"86"),
   142 => (x"d4",x"ff",x"87",x"ca"),
   143 => (x"78",x"ff",x"c3",x"48"),
   144 => (x"87",x"cb",x"48",x"c1"),
   145 => (x"c1",x"87",x"f1",x"fd"),
   146 => (x"db",x"ff",x"05",x"8b"),
   147 => (x"fb",x"48",x"c0",x"87"),
   148 => (x"5e",x"0e",x"87",x"f1"),
   149 => (x"ff",x"0e",x"5c",x"5b"),
   150 => (x"db",x"fd",x"4c",x"d4"),
   151 => (x"1e",x"ea",x"c6",x"87"),
   152 => (x"c1",x"f0",x"e1",x"c0"),
   153 => (x"de",x"fb",x"49",x"c8"),
   154 => (x"c1",x"86",x"c4",x"87"),
   155 => (x"87",x"c8",x"02",x"a8"),
   156 => (x"c0",x"87",x"ea",x"fe"),
   157 => (x"87",x"e2",x"c1",x"48"),
   158 => (x"70",x"87",x"da",x"fa"),
   159 => (x"ff",x"ff",x"cf",x"49"),
   160 => (x"a9",x"ea",x"c6",x"99"),
   161 => (x"fe",x"87",x"c8",x"02"),
   162 => (x"48",x"c0",x"87",x"d3"),
   163 => (x"c3",x"87",x"cb",x"c1"),
   164 => (x"f1",x"c0",x"7c",x"ff"),
   165 => (x"87",x"f4",x"fc",x"4b"),
   166 => (x"c0",x"02",x"98",x"70"),
   167 => (x"1e",x"c0",x"87",x"eb"),
   168 => (x"c1",x"f0",x"ff",x"c0"),
   169 => (x"de",x"fa",x"49",x"fa"),
   170 => (x"70",x"86",x"c4",x"87"),
   171 => (x"87",x"d9",x"05",x"98"),
   172 => (x"6c",x"7c",x"ff",x"c3"),
   173 => (x"7c",x"ff",x"c3",x"49"),
   174 => (x"c1",x"7c",x"7c",x"7c"),
   175 => (x"c4",x"02",x"99",x"c0"),
   176 => (x"d5",x"48",x"c1",x"87"),
   177 => (x"d1",x"48",x"c0",x"87"),
   178 => (x"05",x"ab",x"c2",x"87"),
   179 => (x"48",x"c0",x"87",x"c4"),
   180 => (x"8b",x"c1",x"87",x"c8"),
   181 => (x"87",x"fd",x"fe",x"05"),
   182 => (x"e4",x"f9",x"48",x"c0"),
   183 => (x"1e",x"73",x"1e",x"87"),
   184 => (x"48",x"fc",x"de",x"c2"),
   185 => (x"4b",x"c7",x"78",x"c1"),
   186 => (x"c2",x"48",x"d0",x"ff"),
   187 => (x"87",x"c8",x"fb",x"78"),
   188 => (x"c3",x"48",x"d0",x"ff"),
   189 => (x"c0",x"1e",x"c0",x"78"),
   190 => (x"c0",x"c1",x"d0",x"e5"),
   191 => (x"87",x"c7",x"f9",x"49"),
   192 => (x"a8",x"c1",x"86",x"c4"),
   193 => (x"4b",x"87",x"c1",x"05"),
   194 => (x"c5",x"05",x"ab",x"c2"),
   195 => (x"c0",x"48",x"c0",x"87"),
   196 => (x"8b",x"c1",x"87",x"f9"),
   197 => (x"87",x"d0",x"ff",x"05"),
   198 => (x"c2",x"87",x"f7",x"fc"),
   199 => (x"70",x"58",x"c0",x"df"),
   200 => (x"87",x"cd",x"05",x"98"),
   201 => (x"ff",x"c0",x"1e",x"c1"),
   202 => (x"49",x"d0",x"c1",x"f0"),
   203 => (x"c4",x"87",x"d8",x"f8"),
   204 => (x"48",x"d4",x"ff",x"86"),
   205 => (x"c4",x"78",x"ff",x"c3"),
   206 => (x"df",x"c2",x"87",x"de"),
   207 => (x"d0",x"ff",x"58",x"c4"),
   208 => (x"ff",x"78",x"c2",x"48"),
   209 => (x"ff",x"c3",x"48",x"d4"),
   210 => (x"f7",x"48",x"c1",x"78"),
   211 => (x"5e",x"0e",x"87",x"f5"),
   212 => (x"0e",x"5d",x"5c",x"5b"),
   213 => (x"ff",x"c3",x"4a",x"71"),
   214 => (x"4c",x"d4",x"ff",x"4d"),
   215 => (x"d0",x"ff",x"7c",x"75"),
   216 => (x"78",x"c3",x"c4",x"48"),
   217 => (x"1e",x"72",x"7c",x"75"),
   218 => (x"c1",x"f0",x"ff",x"c0"),
   219 => (x"d6",x"f7",x"49",x"d8"),
   220 => (x"70",x"86",x"c4",x"87"),
   221 => (x"87",x"c5",x"02",x"98"),
   222 => (x"f0",x"c0",x"48",x"c1"),
   223 => (x"c3",x"7c",x"75",x"87"),
   224 => (x"c0",x"c8",x"7c",x"fe"),
   225 => (x"49",x"66",x"d4",x"1e"),
   226 => (x"c4",x"87",x"fa",x"f4"),
   227 => (x"75",x"7c",x"75",x"86"),
   228 => (x"d8",x"7c",x"75",x"7c"),
   229 => (x"75",x"4b",x"e0",x"da"),
   230 => (x"99",x"49",x"6c",x"7c"),
   231 => (x"c1",x"87",x"c5",x"05"),
   232 => (x"87",x"f3",x"05",x"8b"),
   233 => (x"d0",x"ff",x"7c",x"75"),
   234 => (x"c0",x"78",x"c2",x"48"),
   235 => (x"87",x"cf",x"f6",x"48"),
   236 => (x"5c",x"5b",x"5e",x"0e"),
   237 => (x"4b",x"71",x"0e",x"5d"),
   238 => (x"ee",x"c5",x"4c",x"c0"),
   239 => (x"ff",x"4a",x"df",x"cd"),
   240 => (x"ff",x"c3",x"48",x"d4"),
   241 => (x"c3",x"49",x"68",x"78"),
   242 => (x"c0",x"05",x"a9",x"fe"),
   243 => (x"4d",x"70",x"87",x"fd"),
   244 => (x"cc",x"02",x"9b",x"73"),
   245 => (x"1e",x"66",x"d0",x"87"),
   246 => (x"cf",x"f4",x"49",x"73"),
   247 => (x"d6",x"86",x"c4",x"87"),
   248 => (x"48",x"d0",x"ff",x"87"),
   249 => (x"c3",x"78",x"d1",x"c4"),
   250 => (x"66",x"d0",x"7d",x"ff"),
   251 => (x"d4",x"88",x"c1",x"48"),
   252 => (x"98",x"70",x"58",x"a6"),
   253 => (x"ff",x"87",x"f0",x"05"),
   254 => (x"ff",x"c3",x"48",x"d4"),
   255 => (x"9b",x"73",x"78",x"78"),
   256 => (x"ff",x"87",x"c5",x"05"),
   257 => (x"78",x"d0",x"48",x"d0"),
   258 => (x"c1",x"4c",x"4a",x"c1"),
   259 => (x"ee",x"fe",x"05",x"8a"),
   260 => (x"f4",x"48",x"74",x"87"),
   261 => (x"73",x"1e",x"87",x"e9"),
   262 => (x"c0",x"4a",x"71",x"1e"),
   263 => (x"48",x"d4",x"ff",x"4b"),
   264 => (x"ff",x"78",x"ff",x"c3"),
   265 => (x"c3",x"c4",x"48",x"d0"),
   266 => (x"48",x"d4",x"ff",x"78"),
   267 => (x"72",x"78",x"ff",x"c3"),
   268 => (x"f0",x"ff",x"c0",x"1e"),
   269 => (x"f4",x"49",x"d1",x"c1"),
   270 => (x"86",x"c4",x"87",x"cd"),
   271 => (x"d2",x"05",x"98",x"70"),
   272 => (x"1e",x"c0",x"c8",x"87"),
   273 => (x"fd",x"49",x"66",x"cc"),
   274 => (x"86",x"c4",x"87",x"e6"),
   275 => (x"d0",x"ff",x"4b",x"70"),
   276 => (x"73",x"78",x"c2",x"48"),
   277 => (x"87",x"eb",x"f3",x"48"),
   278 => (x"5c",x"5b",x"5e",x"0e"),
   279 => (x"1e",x"c0",x"0e",x"5d"),
   280 => (x"c1",x"f0",x"ff",x"c0"),
   281 => (x"de",x"f3",x"49",x"c9"),
   282 => (x"c2",x"1e",x"d2",x"87"),
   283 => (x"fc",x"49",x"c4",x"df"),
   284 => (x"86",x"c8",x"87",x"fe"),
   285 => (x"84",x"c1",x"4c",x"c0"),
   286 => (x"04",x"ac",x"b7",x"d2"),
   287 => (x"df",x"c2",x"87",x"f8"),
   288 => (x"49",x"bf",x"97",x"c4"),
   289 => (x"c1",x"99",x"c0",x"c3"),
   290 => (x"c0",x"05",x"a9",x"c0"),
   291 => (x"df",x"c2",x"87",x"e7"),
   292 => (x"49",x"bf",x"97",x"cb"),
   293 => (x"df",x"c2",x"31",x"d0"),
   294 => (x"4a",x"bf",x"97",x"cc"),
   295 => (x"b1",x"72",x"32",x"c8"),
   296 => (x"97",x"cd",x"df",x"c2"),
   297 => (x"71",x"b1",x"4a",x"bf"),
   298 => (x"ff",x"ff",x"cf",x"4c"),
   299 => (x"84",x"c1",x"9c",x"ff"),
   300 => (x"e7",x"c1",x"34",x"ca"),
   301 => (x"cd",x"df",x"c2",x"87"),
   302 => (x"c1",x"49",x"bf",x"97"),
   303 => (x"c2",x"99",x"c6",x"31"),
   304 => (x"bf",x"97",x"ce",x"df"),
   305 => (x"2a",x"b7",x"c7",x"4a"),
   306 => (x"df",x"c2",x"b1",x"72"),
   307 => (x"4a",x"bf",x"97",x"c9"),
   308 => (x"c2",x"9d",x"cf",x"4d"),
   309 => (x"bf",x"97",x"ca",x"df"),
   310 => (x"ca",x"9a",x"c3",x"4a"),
   311 => (x"cb",x"df",x"c2",x"32"),
   312 => (x"c2",x"4b",x"bf",x"97"),
   313 => (x"c2",x"b2",x"73",x"33"),
   314 => (x"bf",x"97",x"cc",x"df"),
   315 => (x"9b",x"c0",x"c3",x"4b"),
   316 => (x"73",x"2b",x"b7",x"c6"),
   317 => (x"c1",x"81",x"c2",x"b2"),
   318 => (x"70",x"30",x"71",x"48"),
   319 => (x"75",x"48",x"c1",x"49"),
   320 => (x"72",x"4d",x"70",x"30"),
   321 => (x"71",x"84",x"c1",x"4c"),
   322 => (x"b7",x"c0",x"c8",x"94"),
   323 => (x"87",x"cc",x"06",x"ad"),
   324 => (x"2d",x"b7",x"34",x"c1"),
   325 => (x"ad",x"b7",x"c0",x"c8"),
   326 => (x"87",x"f4",x"ff",x"01"),
   327 => (x"de",x"f0",x"48",x"74"),
   328 => (x"5b",x"5e",x"0e",x"87"),
   329 => (x"f8",x"0e",x"5d",x"5c"),
   330 => (x"ea",x"e7",x"c2",x"86"),
   331 => (x"c2",x"78",x"c0",x"48"),
   332 => (x"c0",x"1e",x"e2",x"df"),
   333 => (x"87",x"de",x"fb",x"49"),
   334 => (x"98",x"70",x"86",x"c4"),
   335 => (x"c0",x"87",x"c5",x"05"),
   336 => (x"87",x"ce",x"c9",x"48"),
   337 => (x"7e",x"c1",x"4d",x"c0"),
   338 => (x"bf",x"c0",x"f3",x"c0"),
   339 => (x"d8",x"e0",x"c2",x"49"),
   340 => (x"4b",x"c8",x"71",x"4a"),
   341 => (x"70",x"87",x"d3",x"ec"),
   342 => (x"87",x"c2",x"05",x"98"),
   343 => (x"f2",x"c0",x"7e",x"c0"),
   344 => (x"c2",x"49",x"bf",x"fc"),
   345 => (x"71",x"4a",x"f4",x"e0"),
   346 => (x"fd",x"eb",x"4b",x"c8"),
   347 => (x"05",x"98",x"70",x"87"),
   348 => (x"7e",x"c0",x"87",x"c2"),
   349 => (x"fd",x"c0",x"02",x"6e"),
   350 => (x"e8",x"e6",x"c2",x"87"),
   351 => (x"e7",x"c2",x"4d",x"bf"),
   352 => (x"7e",x"bf",x"9f",x"e0"),
   353 => (x"ea",x"d6",x"c5",x"48"),
   354 => (x"87",x"c7",x"05",x"a8"),
   355 => (x"bf",x"e8",x"e6",x"c2"),
   356 => (x"6e",x"87",x"ce",x"4d"),
   357 => (x"d5",x"e9",x"ca",x"48"),
   358 => (x"87",x"c5",x"02",x"a8"),
   359 => (x"f1",x"c7",x"48",x"c0"),
   360 => (x"e2",x"df",x"c2",x"87"),
   361 => (x"f9",x"49",x"75",x"1e"),
   362 => (x"86",x"c4",x"87",x"ec"),
   363 => (x"c5",x"05",x"98",x"70"),
   364 => (x"c7",x"48",x"c0",x"87"),
   365 => (x"f2",x"c0",x"87",x"dc"),
   366 => (x"c2",x"49",x"bf",x"fc"),
   367 => (x"71",x"4a",x"f4",x"e0"),
   368 => (x"e5",x"ea",x"4b",x"c8"),
   369 => (x"05",x"98",x"70",x"87"),
   370 => (x"e7",x"c2",x"87",x"c8"),
   371 => (x"78",x"c1",x"48",x"ea"),
   372 => (x"f3",x"c0",x"87",x"da"),
   373 => (x"c2",x"49",x"bf",x"c0"),
   374 => (x"71",x"4a",x"d8",x"e0"),
   375 => (x"c9",x"ea",x"4b",x"c8"),
   376 => (x"02",x"98",x"70",x"87"),
   377 => (x"c0",x"87",x"c5",x"c0"),
   378 => (x"87",x"e6",x"c6",x"48"),
   379 => (x"97",x"e0",x"e7",x"c2"),
   380 => (x"d5",x"c1",x"49",x"bf"),
   381 => (x"cd",x"c0",x"05",x"a9"),
   382 => (x"e1",x"e7",x"c2",x"87"),
   383 => (x"c2",x"49",x"bf",x"97"),
   384 => (x"c0",x"02",x"a9",x"ea"),
   385 => (x"48",x"c0",x"87",x"c5"),
   386 => (x"c2",x"87",x"c7",x"c6"),
   387 => (x"bf",x"97",x"e2",x"df"),
   388 => (x"e9",x"c3",x"48",x"7e"),
   389 => (x"ce",x"c0",x"02",x"a8"),
   390 => (x"c3",x"48",x"6e",x"87"),
   391 => (x"c0",x"02",x"a8",x"eb"),
   392 => (x"48",x"c0",x"87",x"c5"),
   393 => (x"c2",x"87",x"eb",x"c5"),
   394 => (x"bf",x"97",x"ed",x"df"),
   395 => (x"c0",x"05",x"99",x"49"),
   396 => (x"df",x"c2",x"87",x"cc"),
   397 => (x"49",x"bf",x"97",x"ee"),
   398 => (x"c0",x"02",x"a9",x"c2"),
   399 => (x"48",x"c0",x"87",x"c5"),
   400 => (x"c2",x"87",x"cf",x"c5"),
   401 => (x"bf",x"97",x"ef",x"df"),
   402 => (x"e6",x"e7",x"c2",x"48"),
   403 => (x"48",x"4c",x"70",x"58"),
   404 => (x"e7",x"c2",x"88",x"c1"),
   405 => (x"df",x"c2",x"58",x"ea"),
   406 => (x"49",x"bf",x"97",x"f0"),
   407 => (x"df",x"c2",x"81",x"75"),
   408 => (x"4a",x"bf",x"97",x"f1"),
   409 => (x"a1",x"72",x"32",x"c8"),
   410 => (x"f7",x"eb",x"c2",x"7e"),
   411 => (x"c2",x"78",x"6e",x"48"),
   412 => (x"bf",x"97",x"f2",x"df"),
   413 => (x"58",x"a6",x"c8",x"48"),
   414 => (x"bf",x"ea",x"e7",x"c2"),
   415 => (x"87",x"d4",x"c2",x"02"),
   416 => (x"bf",x"fc",x"f2",x"c0"),
   417 => (x"f4",x"e0",x"c2",x"49"),
   418 => (x"4b",x"c8",x"71",x"4a"),
   419 => (x"70",x"87",x"db",x"e7"),
   420 => (x"c5",x"c0",x"02",x"98"),
   421 => (x"c3",x"48",x"c0",x"87"),
   422 => (x"e7",x"c2",x"87",x"f8"),
   423 => (x"c2",x"4c",x"bf",x"e2"),
   424 => (x"c2",x"5c",x"cb",x"ec"),
   425 => (x"bf",x"97",x"c7",x"e0"),
   426 => (x"c2",x"31",x"c8",x"49"),
   427 => (x"bf",x"97",x"c6",x"e0"),
   428 => (x"c2",x"49",x"a1",x"4a"),
   429 => (x"bf",x"97",x"c8",x"e0"),
   430 => (x"72",x"32",x"d0",x"4a"),
   431 => (x"e0",x"c2",x"49",x"a1"),
   432 => (x"4a",x"bf",x"97",x"c9"),
   433 => (x"a1",x"72",x"32",x"d8"),
   434 => (x"91",x"66",x"c4",x"49"),
   435 => (x"bf",x"f7",x"eb",x"c2"),
   436 => (x"ff",x"eb",x"c2",x"81"),
   437 => (x"cf",x"e0",x"c2",x"59"),
   438 => (x"c8",x"4a",x"bf",x"97"),
   439 => (x"ce",x"e0",x"c2",x"32"),
   440 => (x"a2",x"4b",x"bf",x"97"),
   441 => (x"d0",x"e0",x"c2",x"4a"),
   442 => (x"d0",x"4b",x"bf",x"97"),
   443 => (x"4a",x"a2",x"73",x"33"),
   444 => (x"97",x"d1",x"e0",x"c2"),
   445 => (x"9b",x"cf",x"4b",x"bf"),
   446 => (x"a2",x"73",x"33",x"d8"),
   447 => (x"c3",x"ec",x"c2",x"4a"),
   448 => (x"ff",x"eb",x"c2",x"5a"),
   449 => (x"8a",x"c2",x"4a",x"bf"),
   450 => (x"ec",x"c2",x"92",x"74"),
   451 => (x"a1",x"72",x"48",x"c3"),
   452 => (x"87",x"ca",x"c1",x"78"),
   453 => (x"97",x"f4",x"df",x"c2"),
   454 => (x"31",x"c8",x"49",x"bf"),
   455 => (x"97",x"f3",x"df",x"c2"),
   456 => (x"49",x"a1",x"4a",x"bf"),
   457 => (x"59",x"f2",x"e7",x"c2"),
   458 => (x"bf",x"ee",x"e7",x"c2"),
   459 => (x"c7",x"31",x"c5",x"49"),
   460 => (x"29",x"c9",x"81",x"ff"),
   461 => (x"59",x"cb",x"ec",x"c2"),
   462 => (x"97",x"f9",x"df",x"c2"),
   463 => (x"32",x"c8",x"4a",x"bf"),
   464 => (x"97",x"f8",x"df",x"c2"),
   465 => (x"4a",x"a2",x"4b",x"bf"),
   466 => (x"6e",x"92",x"66",x"c4"),
   467 => (x"c7",x"ec",x"c2",x"82"),
   468 => (x"ff",x"eb",x"c2",x"5a"),
   469 => (x"c2",x"78",x"c0",x"48"),
   470 => (x"72",x"48",x"fb",x"eb"),
   471 => (x"ec",x"c2",x"78",x"a1"),
   472 => (x"eb",x"c2",x"48",x"cb"),
   473 => (x"c2",x"78",x"bf",x"ff"),
   474 => (x"c2",x"48",x"cf",x"ec"),
   475 => (x"78",x"bf",x"c3",x"ec"),
   476 => (x"bf",x"ea",x"e7",x"c2"),
   477 => (x"87",x"c9",x"c0",x"02"),
   478 => (x"30",x"c4",x"48",x"74"),
   479 => (x"c9",x"c0",x"7e",x"70"),
   480 => (x"c7",x"ec",x"c2",x"87"),
   481 => (x"30",x"c4",x"48",x"bf"),
   482 => (x"e7",x"c2",x"7e",x"70"),
   483 => (x"78",x"6e",x"48",x"ee"),
   484 => (x"8e",x"f8",x"48",x"c1"),
   485 => (x"4c",x"26",x"4d",x"26"),
   486 => (x"4f",x"26",x"4b",x"26"),
   487 => (x"5c",x"5b",x"5e",x"0e"),
   488 => (x"4a",x"71",x"0e",x"5d"),
   489 => (x"bf",x"ea",x"e7",x"c2"),
   490 => (x"72",x"87",x"cb",x"02"),
   491 => (x"72",x"2b",x"c7",x"4b"),
   492 => (x"9c",x"ff",x"c1",x"4c"),
   493 => (x"4b",x"72",x"87",x"c9"),
   494 => (x"4c",x"72",x"2b",x"c8"),
   495 => (x"c2",x"9c",x"ff",x"c3"),
   496 => (x"83",x"bf",x"f7",x"eb"),
   497 => (x"bf",x"f8",x"f2",x"c0"),
   498 => (x"87",x"d9",x"02",x"ab"),
   499 => (x"5b",x"fc",x"f2",x"c0"),
   500 => (x"1e",x"e2",x"df",x"c2"),
   501 => (x"fd",x"f0",x"49",x"73"),
   502 => (x"70",x"86",x"c4",x"87"),
   503 => (x"87",x"c5",x"05",x"98"),
   504 => (x"e6",x"c0",x"48",x"c0"),
   505 => (x"ea",x"e7",x"c2",x"87"),
   506 => (x"87",x"d2",x"02",x"bf"),
   507 => (x"91",x"c4",x"49",x"74"),
   508 => (x"81",x"e2",x"df",x"c2"),
   509 => (x"ff",x"cf",x"4d",x"69"),
   510 => (x"9d",x"ff",x"ff",x"ff"),
   511 => (x"49",x"74",x"87",x"cb"),
   512 => (x"df",x"c2",x"91",x"c2"),
   513 => (x"69",x"9f",x"81",x"e2"),
   514 => (x"fe",x"48",x"75",x"4d"),
   515 => (x"5e",x"0e",x"87",x"c6"),
   516 => (x"0e",x"5d",x"5c",x"5b"),
   517 => (x"c0",x"4d",x"71",x"1e"),
   518 => (x"ca",x"49",x"c1",x"1e"),
   519 => (x"86",x"c4",x"87",x"ff"),
   520 => (x"02",x"9c",x"4c",x"70"),
   521 => (x"c2",x"87",x"c0",x"c1"),
   522 => (x"75",x"4a",x"f2",x"e7"),
   523 => (x"87",x"df",x"e0",x"49"),
   524 => (x"c0",x"02",x"98",x"70"),
   525 => (x"4a",x"74",x"87",x"f1"),
   526 => (x"4b",x"cb",x"49",x"75"),
   527 => (x"70",x"87",x"c5",x"e1"),
   528 => (x"e2",x"c0",x"02",x"98"),
   529 => (x"74",x"1e",x"c0",x"87"),
   530 => (x"87",x"c7",x"02",x"9c"),
   531 => (x"c0",x"48",x"a6",x"c4"),
   532 => (x"c4",x"87",x"c5",x"78"),
   533 => (x"78",x"c1",x"48",x"a6"),
   534 => (x"c9",x"49",x"66",x"c4"),
   535 => (x"86",x"c4",x"87",x"ff"),
   536 => (x"05",x"9c",x"4c",x"70"),
   537 => (x"74",x"87",x"c0",x"ff"),
   538 => (x"e7",x"fc",x"26",x"48"),
   539 => (x"5b",x"5e",x"0e",x"87"),
   540 => (x"1e",x"0e",x"5d",x"5c"),
   541 => (x"05",x"9b",x"4b",x"71"),
   542 => (x"48",x"c0",x"87",x"c5"),
   543 => (x"c8",x"87",x"e5",x"c1"),
   544 => (x"7d",x"c0",x"4d",x"a3"),
   545 => (x"c7",x"02",x"66",x"d4"),
   546 => (x"97",x"66",x"d4",x"87"),
   547 => (x"87",x"c5",x"05",x"bf"),
   548 => (x"cf",x"c1",x"48",x"c0"),
   549 => (x"49",x"66",x"d4",x"87"),
   550 => (x"70",x"87",x"f3",x"fd"),
   551 => (x"c1",x"02",x"9c",x"4c"),
   552 => (x"a4",x"dc",x"87",x"c0"),
   553 => (x"da",x"7d",x"69",x"49"),
   554 => (x"a3",x"c4",x"49",x"a4"),
   555 => (x"7a",x"69",x"9f",x"4a"),
   556 => (x"bf",x"ea",x"e7",x"c2"),
   557 => (x"d4",x"87",x"d2",x"02"),
   558 => (x"69",x"9f",x"49",x"a4"),
   559 => (x"ff",x"ff",x"c0",x"49"),
   560 => (x"d0",x"48",x"71",x"99"),
   561 => (x"c2",x"7e",x"70",x"30"),
   562 => (x"6e",x"7e",x"c0",x"87"),
   563 => (x"80",x"6a",x"48",x"49"),
   564 => (x"7b",x"c0",x"7a",x"70"),
   565 => (x"6a",x"49",x"a3",x"cc"),
   566 => (x"49",x"a3",x"d0",x"79"),
   567 => (x"48",x"c1",x"79",x"c0"),
   568 => (x"48",x"c0",x"87",x"c2"),
   569 => (x"87",x"ec",x"fa",x"26"),
   570 => (x"5c",x"5b",x"5e",x"0e"),
   571 => (x"4c",x"71",x"0e",x"5d"),
   572 => (x"ca",x"c1",x"02",x"9c"),
   573 => (x"49",x"a4",x"c8",x"87"),
   574 => (x"c2",x"c1",x"02",x"69"),
   575 => (x"4a",x"66",x"d0",x"87"),
   576 => (x"d4",x"82",x"49",x"6c"),
   577 => (x"66",x"d0",x"5a",x"a6"),
   578 => (x"e7",x"c2",x"b9",x"4d"),
   579 => (x"ff",x"4a",x"bf",x"e6"),
   580 => (x"71",x"99",x"72",x"ba"),
   581 => (x"e4",x"c0",x"02",x"99"),
   582 => (x"4b",x"a4",x"c4",x"87"),
   583 => (x"fb",x"f9",x"49",x"6b"),
   584 => (x"c2",x"7b",x"70",x"87"),
   585 => (x"49",x"bf",x"e2",x"e7"),
   586 => (x"7c",x"71",x"81",x"6c"),
   587 => (x"e7",x"c2",x"b9",x"75"),
   588 => (x"ff",x"4a",x"bf",x"e6"),
   589 => (x"71",x"99",x"72",x"ba"),
   590 => (x"dc",x"ff",x"05",x"99"),
   591 => (x"f9",x"7c",x"75",x"87"),
   592 => (x"73",x"1e",x"87",x"d2"),
   593 => (x"9b",x"4b",x"71",x"1e"),
   594 => (x"c8",x"87",x"c7",x"02"),
   595 => (x"05",x"69",x"49",x"a3"),
   596 => (x"48",x"c0",x"87",x"c5"),
   597 => (x"c2",x"87",x"f7",x"c0"),
   598 => (x"4a",x"bf",x"fb",x"eb"),
   599 => (x"69",x"49",x"a3",x"c4"),
   600 => (x"c2",x"89",x"c2",x"49"),
   601 => (x"91",x"bf",x"e2",x"e7"),
   602 => (x"c2",x"4a",x"a2",x"71"),
   603 => (x"49",x"bf",x"e6",x"e7"),
   604 => (x"a2",x"71",x"99",x"6b"),
   605 => (x"fc",x"f2",x"c0",x"4a"),
   606 => (x"1e",x"66",x"c8",x"5a"),
   607 => (x"d5",x"ea",x"49",x"72"),
   608 => (x"70",x"86",x"c4",x"87"),
   609 => (x"87",x"c4",x"05",x"98"),
   610 => (x"87",x"c2",x"48",x"c0"),
   611 => (x"c7",x"f8",x"48",x"c1"),
   612 => (x"1e",x"73",x"1e",x"87"),
   613 => (x"02",x"9b",x"4b",x"71"),
   614 => (x"a3",x"c8",x"87",x"c7"),
   615 => (x"c5",x"05",x"69",x"49"),
   616 => (x"c0",x"48",x"c0",x"87"),
   617 => (x"eb",x"c2",x"87",x"f7"),
   618 => (x"c4",x"4a",x"bf",x"fb"),
   619 => (x"49",x"69",x"49",x"a3"),
   620 => (x"e7",x"c2",x"89",x"c2"),
   621 => (x"71",x"91",x"bf",x"e2"),
   622 => (x"e7",x"c2",x"4a",x"a2"),
   623 => (x"6b",x"49",x"bf",x"e6"),
   624 => (x"4a",x"a2",x"71",x"99"),
   625 => (x"5a",x"fc",x"f2",x"c0"),
   626 => (x"72",x"1e",x"66",x"c8"),
   627 => (x"87",x"fe",x"e5",x"49"),
   628 => (x"98",x"70",x"86",x"c4"),
   629 => (x"c0",x"87",x"c4",x"05"),
   630 => (x"c1",x"87",x"c2",x"48"),
   631 => (x"87",x"f8",x"f6",x"48"),
   632 => (x"5c",x"5b",x"5e",x"0e"),
   633 => (x"71",x"1e",x"0e",x"5d"),
   634 => (x"4c",x"66",x"d4",x"4b"),
   635 => (x"9b",x"73",x"2c",x"c9"),
   636 => (x"87",x"cf",x"c1",x"02"),
   637 => (x"69",x"49",x"a3",x"c8"),
   638 => (x"87",x"c7",x"c1",x"02"),
   639 => (x"d4",x"4d",x"a3",x"d0"),
   640 => (x"e7",x"c2",x"7d",x"66"),
   641 => (x"ff",x"49",x"bf",x"e6"),
   642 => (x"99",x"4a",x"6b",x"b9"),
   643 => (x"03",x"ac",x"71",x"7e"),
   644 => (x"7b",x"c0",x"87",x"cd"),
   645 => (x"4a",x"a3",x"cc",x"7d"),
   646 => (x"6a",x"49",x"a3",x"c4"),
   647 => (x"72",x"87",x"c2",x"79"),
   648 => (x"02",x"9c",x"74",x"8c"),
   649 => (x"1e",x"49",x"87",x"dd"),
   650 => (x"fb",x"fa",x"49",x"73"),
   651 => (x"d4",x"86",x"c4",x"87"),
   652 => (x"ff",x"c7",x"49",x"66"),
   653 => (x"87",x"cb",x"02",x"99"),
   654 => (x"1e",x"e2",x"df",x"c2"),
   655 => (x"c1",x"fc",x"49",x"73"),
   656 => (x"26",x"86",x"c4",x"87"),
   657 => (x"1e",x"87",x"cd",x"f5"),
   658 => (x"4b",x"71",x"1e",x"73"),
   659 => (x"e4",x"c0",x"02",x"9b"),
   660 => (x"cf",x"ec",x"c2",x"87"),
   661 => (x"c2",x"4a",x"73",x"5b"),
   662 => (x"e2",x"e7",x"c2",x"8a"),
   663 => (x"c2",x"92",x"49",x"bf"),
   664 => (x"48",x"bf",x"fb",x"eb"),
   665 => (x"ec",x"c2",x"80",x"72"),
   666 => (x"48",x"71",x"58",x"d3"),
   667 => (x"e7",x"c2",x"30",x"c4"),
   668 => (x"ed",x"c0",x"58",x"f2"),
   669 => (x"cb",x"ec",x"c2",x"87"),
   670 => (x"ff",x"eb",x"c2",x"48"),
   671 => (x"ec",x"c2",x"78",x"bf"),
   672 => (x"ec",x"c2",x"48",x"cf"),
   673 => (x"c2",x"78",x"bf",x"c3"),
   674 => (x"02",x"bf",x"ea",x"e7"),
   675 => (x"e7",x"c2",x"87",x"c9"),
   676 => (x"c4",x"49",x"bf",x"e2"),
   677 => (x"c2",x"87",x"c7",x"31"),
   678 => (x"49",x"bf",x"c7",x"ec"),
   679 => (x"e7",x"c2",x"31",x"c4"),
   680 => (x"f3",x"f3",x"59",x"f2"),
   681 => (x"5b",x"5e",x"0e",x"87"),
   682 => (x"4a",x"71",x"0e",x"5c"),
   683 => (x"9a",x"72",x"4b",x"c0"),
   684 => (x"87",x"e1",x"c0",x"02"),
   685 => (x"9f",x"49",x"a2",x"da"),
   686 => (x"e7",x"c2",x"4b",x"69"),
   687 => (x"cf",x"02",x"bf",x"ea"),
   688 => (x"49",x"a2",x"d4",x"87"),
   689 => (x"4c",x"49",x"69",x"9f"),
   690 => (x"9c",x"ff",x"ff",x"c0"),
   691 => (x"87",x"c2",x"34",x"d0"),
   692 => (x"49",x"74",x"4c",x"c0"),
   693 => (x"fd",x"49",x"73",x"b3"),
   694 => (x"f9",x"f2",x"87",x"ed"),
   695 => (x"5b",x"5e",x"0e",x"87"),
   696 => (x"f4",x"0e",x"5d",x"5c"),
   697 => (x"c0",x"4a",x"71",x"86"),
   698 => (x"02",x"9a",x"72",x"7e"),
   699 => (x"df",x"c2",x"87",x"d8"),
   700 => (x"78",x"c0",x"48",x"de"),
   701 => (x"48",x"d6",x"df",x"c2"),
   702 => (x"bf",x"cf",x"ec",x"c2"),
   703 => (x"da",x"df",x"c2",x"78"),
   704 => (x"cb",x"ec",x"c2",x"48"),
   705 => (x"e7",x"c2",x"78",x"bf"),
   706 => (x"50",x"c0",x"48",x"ff"),
   707 => (x"bf",x"ee",x"e7",x"c2"),
   708 => (x"de",x"df",x"c2",x"49"),
   709 => (x"aa",x"71",x"4a",x"bf"),
   710 => (x"87",x"c9",x"c4",x"03"),
   711 => (x"99",x"cf",x"49",x"72"),
   712 => (x"87",x"e9",x"c0",x"05"),
   713 => (x"48",x"f8",x"f2",x"c0"),
   714 => (x"bf",x"d6",x"df",x"c2"),
   715 => (x"e2",x"df",x"c2",x"78"),
   716 => (x"d6",x"df",x"c2",x"1e"),
   717 => (x"df",x"c2",x"49",x"bf"),
   718 => (x"a1",x"c1",x"48",x"d6"),
   719 => (x"d5",x"e3",x"71",x"78"),
   720 => (x"c0",x"86",x"c4",x"87"),
   721 => (x"c2",x"48",x"f4",x"f2"),
   722 => (x"cc",x"78",x"e2",x"df"),
   723 => (x"f4",x"f2",x"c0",x"87"),
   724 => (x"e0",x"c0",x"48",x"bf"),
   725 => (x"f8",x"f2",x"c0",x"80"),
   726 => (x"de",x"df",x"c2",x"58"),
   727 => (x"80",x"c1",x"48",x"bf"),
   728 => (x"58",x"e2",x"df",x"c2"),
   729 => (x"00",x"0c",x"b4",x"27"),
   730 => (x"bf",x"97",x"bf",x"00"),
   731 => (x"c2",x"02",x"9d",x"4d"),
   732 => (x"e5",x"c3",x"87",x"e3"),
   733 => (x"dc",x"c2",x"02",x"ad"),
   734 => (x"f4",x"f2",x"c0",x"87"),
   735 => (x"a3",x"cb",x"4b",x"bf"),
   736 => (x"cf",x"4c",x"11",x"49"),
   737 => (x"d2",x"c1",x"05",x"ac"),
   738 => (x"df",x"49",x"75",x"87"),
   739 => (x"cd",x"89",x"c1",x"99"),
   740 => (x"f2",x"e7",x"c2",x"91"),
   741 => (x"4a",x"a3",x"c1",x"81"),
   742 => (x"a3",x"c3",x"51",x"12"),
   743 => (x"c5",x"51",x"12",x"4a"),
   744 => (x"51",x"12",x"4a",x"a3"),
   745 => (x"12",x"4a",x"a3",x"c7"),
   746 => (x"4a",x"a3",x"c9",x"51"),
   747 => (x"a3",x"ce",x"51",x"12"),
   748 => (x"d0",x"51",x"12",x"4a"),
   749 => (x"51",x"12",x"4a",x"a3"),
   750 => (x"12",x"4a",x"a3",x"d2"),
   751 => (x"4a",x"a3",x"d4",x"51"),
   752 => (x"a3",x"d6",x"51",x"12"),
   753 => (x"d8",x"51",x"12",x"4a"),
   754 => (x"51",x"12",x"4a",x"a3"),
   755 => (x"12",x"4a",x"a3",x"dc"),
   756 => (x"4a",x"a3",x"de",x"51"),
   757 => (x"7e",x"c1",x"51",x"12"),
   758 => (x"74",x"87",x"fa",x"c0"),
   759 => (x"05",x"99",x"c8",x"49"),
   760 => (x"74",x"87",x"eb",x"c0"),
   761 => (x"05",x"99",x"d0",x"49"),
   762 => (x"66",x"dc",x"87",x"d1"),
   763 => (x"87",x"cb",x"c0",x"02"),
   764 => (x"66",x"dc",x"49",x"73"),
   765 => (x"02",x"98",x"70",x"0f"),
   766 => (x"6e",x"87",x"d3",x"c0"),
   767 => (x"87",x"c6",x"c0",x"05"),
   768 => (x"48",x"f2",x"e7",x"c2"),
   769 => (x"f2",x"c0",x"50",x"c0"),
   770 => (x"c2",x"48",x"bf",x"f4"),
   771 => (x"e7",x"c2",x"87",x"e1"),
   772 => (x"50",x"c0",x"48",x"ff"),
   773 => (x"ee",x"e7",x"c2",x"7e"),
   774 => (x"df",x"c2",x"49",x"bf"),
   775 => (x"71",x"4a",x"bf",x"de"),
   776 => (x"f7",x"fb",x"04",x"aa"),
   777 => (x"cf",x"ec",x"c2",x"87"),
   778 => (x"c8",x"c0",x"05",x"bf"),
   779 => (x"ea",x"e7",x"c2",x"87"),
   780 => (x"f8",x"c1",x"02",x"bf"),
   781 => (x"da",x"df",x"c2",x"87"),
   782 => (x"df",x"ed",x"49",x"bf"),
   783 => (x"c2",x"49",x"70",x"87"),
   784 => (x"c4",x"59",x"de",x"df"),
   785 => (x"df",x"c2",x"48",x"a6"),
   786 => (x"c2",x"78",x"bf",x"da"),
   787 => (x"02",x"bf",x"ea",x"e7"),
   788 => (x"c4",x"87",x"d8",x"c0"),
   789 => (x"ff",x"cf",x"49",x"66"),
   790 => (x"99",x"f8",x"ff",x"ff"),
   791 => (x"c5",x"c0",x"02",x"a9"),
   792 => (x"c0",x"4c",x"c0",x"87"),
   793 => (x"4c",x"c1",x"87",x"e1"),
   794 => (x"c4",x"87",x"dc",x"c0"),
   795 => (x"ff",x"cf",x"49",x"66"),
   796 => (x"02",x"a9",x"99",x"f8"),
   797 => (x"c8",x"87",x"c8",x"c0"),
   798 => (x"78",x"c0",x"48",x"a6"),
   799 => (x"c8",x"87",x"c5",x"c0"),
   800 => (x"78",x"c1",x"48",x"a6"),
   801 => (x"74",x"4c",x"66",x"c8"),
   802 => (x"e0",x"c0",x"05",x"9c"),
   803 => (x"49",x"66",x"c4",x"87"),
   804 => (x"e7",x"c2",x"89",x"c2"),
   805 => (x"91",x"4a",x"bf",x"e2"),
   806 => (x"bf",x"fb",x"eb",x"c2"),
   807 => (x"d6",x"df",x"c2",x"4a"),
   808 => (x"78",x"a1",x"72",x"48"),
   809 => (x"48",x"de",x"df",x"c2"),
   810 => (x"df",x"f9",x"78",x"c0"),
   811 => (x"f4",x"48",x"c0",x"87"),
   812 => (x"87",x"e0",x"eb",x"8e"),
   813 => (x"00",x"00",x"00",x"00"),
   814 => (x"ff",x"ff",x"ff",x"ff"),
   815 => (x"00",x"00",x"0c",x"c4"),
   816 => (x"00",x"00",x"0c",x"cd"),
   817 => (x"33",x"54",x"41",x"46"),
   818 => (x"20",x"20",x"20",x"32"),
   819 => (x"54",x"41",x"46",x"00"),
   820 => (x"20",x"20",x"36",x"31"),
   821 => (x"ff",x"1e",x"00",x"20"),
   822 => (x"ff",x"c3",x"48",x"d4"),
   823 => (x"26",x"48",x"68",x"78"),
   824 => (x"d4",x"ff",x"1e",x"4f"),
   825 => (x"78",x"ff",x"c3",x"48"),
   826 => (x"c8",x"48",x"d0",x"ff"),
   827 => (x"d4",x"ff",x"78",x"e1"),
   828 => (x"c2",x"78",x"d4",x"48"),
   829 => (x"ff",x"48",x"d3",x"ec"),
   830 => (x"26",x"50",x"bf",x"d4"),
   831 => (x"d0",x"ff",x"1e",x"4f"),
   832 => (x"78",x"e0",x"c0",x"48"),
   833 => (x"ff",x"1e",x"4f",x"26"),
   834 => (x"49",x"70",x"87",x"cc"),
   835 => (x"87",x"c6",x"02",x"99"),
   836 => (x"05",x"a9",x"fb",x"c0"),
   837 => (x"48",x"71",x"87",x"f1"),
   838 => (x"5e",x"0e",x"4f",x"26"),
   839 => (x"71",x"0e",x"5c",x"5b"),
   840 => (x"fe",x"4c",x"c0",x"4b"),
   841 => (x"49",x"70",x"87",x"f0"),
   842 => (x"f9",x"c0",x"02",x"99"),
   843 => (x"a9",x"ec",x"c0",x"87"),
   844 => (x"87",x"f2",x"c0",x"02"),
   845 => (x"02",x"a9",x"fb",x"c0"),
   846 => (x"cc",x"87",x"eb",x"c0"),
   847 => (x"03",x"ac",x"b7",x"66"),
   848 => (x"66",x"d0",x"87",x"c7"),
   849 => (x"71",x"87",x"c2",x"02"),
   850 => (x"02",x"99",x"71",x"53"),
   851 => (x"84",x"c1",x"87",x"c2"),
   852 => (x"70",x"87",x"c3",x"fe"),
   853 => (x"cd",x"02",x"99",x"49"),
   854 => (x"a9",x"ec",x"c0",x"87"),
   855 => (x"c0",x"87",x"c7",x"02"),
   856 => (x"ff",x"05",x"a9",x"fb"),
   857 => (x"66",x"d0",x"87",x"d5"),
   858 => (x"c0",x"87",x"c3",x"02"),
   859 => (x"ec",x"c0",x"7b",x"97"),
   860 => (x"87",x"c4",x"05",x"a9"),
   861 => (x"87",x"c5",x"4a",x"74"),
   862 => (x"0a",x"c0",x"4a",x"74"),
   863 => (x"c2",x"48",x"72",x"8a"),
   864 => (x"26",x"4d",x"26",x"87"),
   865 => (x"26",x"4b",x"26",x"4c"),
   866 => (x"c9",x"fd",x"1e",x"4f"),
   867 => (x"c0",x"49",x"70",x"87"),
   868 => (x"04",x"a9",x"b7",x"f0"),
   869 => (x"f9",x"c0",x"87",x"ca"),
   870 => (x"c3",x"01",x"a9",x"b7"),
   871 => (x"89",x"f0",x"c0",x"87"),
   872 => (x"a9",x"b7",x"c1",x"c1"),
   873 => (x"c1",x"87",x"ca",x"04"),
   874 => (x"01",x"a9",x"b7",x"da"),
   875 => (x"f7",x"c0",x"87",x"c3"),
   876 => (x"b7",x"e1",x"c1",x"89"),
   877 => (x"87",x"ca",x"04",x"a9"),
   878 => (x"a9",x"b7",x"fa",x"c1"),
   879 => (x"c0",x"87",x"c3",x"01"),
   880 => (x"48",x"71",x"89",x"fd"),
   881 => (x"5e",x"0e",x"4f",x"26"),
   882 => (x"71",x"0e",x"5c",x"5b"),
   883 => (x"4c",x"d4",x"ff",x"4a"),
   884 => (x"ea",x"c0",x"49",x"72"),
   885 => (x"9b",x"4b",x"70",x"87"),
   886 => (x"c1",x"87",x"c2",x"02"),
   887 => (x"48",x"d0",x"ff",x"8b"),
   888 => (x"c1",x"78",x"c5",x"c8"),
   889 => (x"49",x"73",x"7c",x"d5"),
   890 => (x"e2",x"c1",x"31",x"c6"),
   891 => (x"4a",x"bf",x"97",x"fe"),
   892 => (x"70",x"b0",x"71",x"48"),
   893 => (x"48",x"d0",x"ff",x"7c"),
   894 => (x"48",x"73",x"78",x"c4"),
   895 => (x"0e",x"87",x"c4",x"fe"),
   896 => (x"5d",x"5c",x"5b",x"5e"),
   897 => (x"71",x"86",x"f8",x"0e"),
   898 => (x"fb",x"7e",x"c0",x"4c"),
   899 => (x"4b",x"c0",x"87",x"d3"),
   900 => (x"97",x"ec",x"fa",x"c0"),
   901 => (x"a9",x"c0",x"49",x"bf"),
   902 => (x"fb",x"87",x"cf",x"04"),
   903 => (x"83",x"c1",x"87",x"e8"),
   904 => (x"97",x"ec",x"fa",x"c0"),
   905 => (x"06",x"ab",x"49",x"bf"),
   906 => (x"fa",x"c0",x"87",x"f1"),
   907 => (x"02",x"bf",x"97",x"ec"),
   908 => (x"e1",x"fa",x"87",x"cf"),
   909 => (x"99",x"49",x"70",x"87"),
   910 => (x"c0",x"87",x"c6",x"02"),
   911 => (x"f1",x"05",x"a9",x"ec"),
   912 => (x"fa",x"4b",x"c0",x"87"),
   913 => (x"4d",x"70",x"87",x"d0"),
   914 => (x"c8",x"87",x"cb",x"fa"),
   915 => (x"c5",x"fa",x"58",x"a6"),
   916 => (x"c1",x"4a",x"70",x"87"),
   917 => (x"49",x"a4",x"c8",x"83"),
   918 => (x"ad",x"49",x"69",x"97"),
   919 => (x"c0",x"87",x"c7",x"02"),
   920 => (x"c0",x"05",x"ad",x"ff"),
   921 => (x"a4",x"c9",x"87",x"e7"),
   922 => (x"49",x"69",x"97",x"49"),
   923 => (x"02",x"a9",x"66",x"c4"),
   924 => (x"c0",x"48",x"87",x"c7"),
   925 => (x"d4",x"05",x"a8",x"ff"),
   926 => (x"49",x"a4",x"ca",x"87"),
   927 => (x"aa",x"49",x"69",x"97"),
   928 => (x"c0",x"87",x"c6",x"02"),
   929 => (x"c4",x"05",x"aa",x"ff"),
   930 => (x"d0",x"7e",x"c1",x"87"),
   931 => (x"ad",x"ec",x"c0",x"87"),
   932 => (x"c0",x"87",x"c6",x"02"),
   933 => (x"c4",x"05",x"ad",x"fb"),
   934 => (x"c1",x"4b",x"c0",x"87"),
   935 => (x"fe",x"02",x"6e",x"7e"),
   936 => (x"d8",x"f9",x"87",x"e1"),
   937 => (x"f8",x"48",x"73",x"87"),
   938 => (x"87",x"d5",x"fb",x"8e"),
   939 => (x"5b",x"5e",x"0e",x"00"),
   940 => (x"1e",x"0e",x"5d",x"5c"),
   941 => (x"d4",x"ff",x"4d",x"71"),
   942 => (x"c2",x"1e",x"75",x"4b"),
   943 => (x"e6",x"49",x"d8",x"ec"),
   944 => (x"86",x"c4",x"87",x"eb"),
   945 => (x"c3",x"02",x"98",x"70"),
   946 => (x"ec",x"c2",x"87",x"d8"),
   947 => (x"75",x"4c",x"bf",x"e0"),
   948 => (x"87",x"f2",x"fb",x"49"),
   949 => (x"c8",x"48",x"d0",x"ff"),
   950 => (x"d6",x"c1",x"78",x"c5"),
   951 => (x"75",x"4a",x"c0",x"7b"),
   952 => (x"7b",x"11",x"49",x"a2"),
   953 => (x"b7",x"cb",x"82",x"c1"),
   954 => (x"87",x"f3",x"04",x"aa"),
   955 => (x"ff",x"c3",x"4a",x"cc"),
   956 => (x"c0",x"82",x"c1",x"7b"),
   957 => (x"04",x"aa",x"b7",x"e0"),
   958 => (x"d0",x"ff",x"87",x"f4"),
   959 => (x"c3",x"78",x"c4",x"48"),
   960 => (x"c5",x"c8",x"7b",x"ff"),
   961 => (x"7b",x"d3",x"c1",x"78"),
   962 => (x"78",x"c4",x"7b",x"c1"),
   963 => (x"c1",x"02",x"9c",x"74"),
   964 => (x"df",x"c2",x"87",x"ff"),
   965 => (x"c0",x"c8",x"7e",x"e2"),
   966 => (x"b7",x"c0",x"8c",x"4d"),
   967 => (x"87",x"c6",x"03",x"ac"),
   968 => (x"4d",x"a4",x"c0",x"c8"),
   969 => (x"c0",x"c8",x"4c",x"c0"),
   970 => (x"87",x"dc",x"05",x"ad"),
   971 => (x"97",x"d3",x"ec",x"c2"),
   972 => (x"99",x"d0",x"49",x"bf"),
   973 => (x"c0",x"87",x"d1",x"02"),
   974 => (x"d8",x"ec",x"c2",x"1e"),
   975 => (x"87",x"c2",x"e8",x"49"),
   976 => (x"49",x"70",x"86",x"c4"),
   977 => (x"87",x"ee",x"c0",x"4a"),
   978 => (x"1e",x"e2",x"df",x"c2"),
   979 => (x"49",x"d8",x"ec",x"c2"),
   980 => (x"c4",x"87",x"ef",x"e7"),
   981 => (x"4a",x"49",x"70",x"86"),
   982 => (x"c8",x"48",x"d0",x"ff"),
   983 => (x"d4",x"c1",x"78",x"c5"),
   984 => (x"bf",x"97",x"6e",x"7b"),
   985 => (x"c1",x"48",x"6e",x"7b"),
   986 => (x"c1",x"7e",x"70",x"80"),
   987 => (x"f0",x"ff",x"05",x"8d"),
   988 => (x"48",x"d0",x"ff",x"87"),
   989 => (x"9a",x"72",x"78",x"c4"),
   990 => (x"c0",x"87",x"c5",x"05"),
   991 => (x"87",x"e4",x"c0",x"48"),
   992 => (x"ec",x"c2",x"1e",x"c1"),
   993 => (x"df",x"e5",x"49",x"d8"),
   994 => (x"74",x"86",x"c4",x"87"),
   995 => (x"c1",x"fe",x"05",x"9c"),
   996 => (x"48",x"d0",x"ff",x"87"),
   997 => (x"c1",x"78",x"c5",x"c8"),
   998 => (x"7b",x"c0",x"7b",x"d3"),
   999 => (x"48",x"c1",x"78",x"c4"),
  1000 => (x"48",x"c0",x"87",x"c2"),
  1001 => (x"26",x"4d",x"26",x"26"),
  1002 => (x"26",x"4b",x"26",x"4c"),
  1003 => (x"5b",x"5e",x"0e",x"4f"),
  1004 => (x"1e",x"0e",x"5d",x"5c"),
  1005 => (x"4c",x"c0",x"4b",x"71"),
  1006 => (x"c0",x"04",x"ab",x"4d"),
  1007 => (x"f7",x"c0",x"87",x"e8"),
  1008 => (x"9d",x"75",x"1e",x"ff"),
  1009 => (x"c0",x"87",x"c4",x"02"),
  1010 => (x"c1",x"87",x"c2",x"4a"),
  1011 => (x"ec",x"49",x"72",x"4a"),
  1012 => (x"86",x"c4",x"87",x"cb"),
  1013 => (x"84",x"c1",x"7e",x"70"),
  1014 => (x"87",x"c2",x"05",x"6e"),
  1015 => (x"85",x"c1",x"4c",x"73"),
  1016 => (x"ff",x"06",x"ac",x"73"),
  1017 => (x"48",x"6e",x"87",x"d8"),
  1018 => (x"87",x"f9",x"fe",x"26"),
  1019 => (x"5c",x"5b",x"5e",x"0e"),
  1020 => (x"cc",x"4b",x"71",x"0e"),
  1021 => (x"87",x"d8",x"02",x"66"),
  1022 => (x"8c",x"f0",x"c0",x"4c"),
  1023 => (x"74",x"87",x"d8",x"02"),
  1024 => (x"02",x"8a",x"c1",x"4a"),
  1025 => (x"02",x"8a",x"87",x"d1"),
  1026 => (x"02",x"8a",x"87",x"cd"),
  1027 => (x"87",x"d9",x"87",x"c9"),
  1028 => (x"d8",x"fa",x"49",x"73"),
  1029 => (x"74",x"87",x"d2",x"87"),
  1030 => (x"c1",x"49",x"c0",x"1e"),
  1031 => (x"74",x"87",x"c8",x"db"),
  1032 => (x"c1",x"49",x"73",x"1e"),
  1033 => (x"c8",x"87",x"c0",x"db"),
  1034 => (x"87",x"fb",x"fd",x"86"),
  1035 => (x"5c",x"5b",x"5e",x"0e"),
  1036 => (x"71",x"1e",x"0e",x"5d"),
  1037 => (x"91",x"de",x"49",x"4c"),
  1038 => (x"4d",x"c0",x"ed",x"c2"),
  1039 => (x"6d",x"97",x"85",x"71"),
  1040 => (x"87",x"dc",x"c1",x"02"),
  1041 => (x"bf",x"ec",x"ec",x"c2"),
  1042 => (x"72",x"82",x"74",x"4a"),
  1043 => (x"87",x"dd",x"fd",x"49"),
  1044 => (x"02",x"6e",x"7e",x"70"),
  1045 => (x"c2",x"87",x"f2",x"c0"),
  1046 => (x"6e",x"4b",x"f4",x"ec"),
  1047 => (x"ff",x"49",x"cb",x"4a"),
  1048 => (x"74",x"87",x"c5",x"c1"),
  1049 => (x"c1",x"93",x"cb",x"4b"),
  1050 => (x"c4",x"83",x"ce",x"e3"),
  1051 => (x"e4",x"c2",x"c1",x"83"),
  1052 => (x"c1",x"49",x"74",x"7b"),
  1053 => (x"75",x"87",x"c0",x"c5"),
  1054 => (x"ff",x"e2",x"c1",x"7b"),
  1055 => (x"1e",x"49",x"bf",x"97"),
  1056 => (x"49",x"f4",x"ec",x"c2"),
  1057 => (x"c4",x"87",x"e5",x"fd"),
  1058 => (x"c1",x"49",x"74",x"86"),
  1059 => (x"c0",x"87",x"e8",x"c4"),
  1060 => (x"c7",x"c6",x"c1",x"49"),
  1061 => (x"d4",x"ec",x"c2",x"87"),
  1062 => (x"c1",x"78",x"c0",x"48"),
  1063 => (x"87",x"ff",x"dc",x"49"),
  1064 => (x"87",x"c1",x"fc",x"26"),
  1065 => (x"64",x"61",x"6f",x"4c"),
  1066 => (x"2e",x"67",x"6e",x"69"),
  1067 => (x"0e",x"00",x"2e",x"2e"),
  1068 => (x"0e",x"5c",x"5b",x"5e"),
  1069 => (x"c2",x"4a",x"4b",x"71"),
  1070 => (x"82",x"bf",x"ec",x"ec"),
  1071 => (x"ec",x"fb",x"49",x"72"),
  1072 => (x"9c",x"4c",x"70",x"87"),
  1073 => (x"49",x"87",x"c4",x"02"),
  1074 => (x"c2",x"87",x"da",x"e7"),
  1075 => (x"c0",x"48",x"ec",x"ec"),
  1076 => (x"dc",x"49",x"c1",x"78"),
  1077 => (x"ce",x"fb",x"87",x"c9"),
  1078 => (x"5b",x"5e",x"0e",x"87"),
  1079 => (x"f4",x"0e",x"5d",x"5c"),
  1080 => (x"e2",x"df",x"c2",x"86"),
  1081 => (x"c4",x"4c",x"c0",x"4d"),
  1082 => (x"78",x"c0",x"48",x"a6"),
  1083 => (x"bf",x"ec",x"ec",x"c2"),
  1084 => (x"06",x"a9",x"c0",x"49"),
  1085 => (x"c2",x"87",x"c1",x"c1"),
  1086 => (x"98",x"48",x"e2",x"df"),
  1087 => (x"87",x"f8",x"c0",x"02"),
  1088 => (x"1e",x"ff",x"f7",x"c0"),
  1089 => (x"c7",x"02",x"66",x"c8"),
  1090 => (x"48",x"a6",x"c4",x"87"),
  1091 => (x"87",x"c5",x"78",x"c0"),
  1092 => (x"c1",x"48",x"a6",x"c4"),
  1093 => (x"49",x"66",x"c4",x"78"),
  1094 => (x"c4",x"87",x"c2",x"e7"),
  1095 => (x"c1",x"4d",x"70",x"86"),
  1096 => (x"48",x"66",x"c4",x"84"),
  1097 => (x"a6",x"c8",x"80",x"c1"),
  1098 => (x"ec",x"ec",x"c2",x"58"),
  1099 => (x"03",x"ac",x"49",x"bf"),
  1100 => (x"9d",x"75",x"87",x"c6"),
  1101 => (x"87",x"c8",x"ff",x"05"),
  1102 => (x"9d",x"75",x"4c",x"c0"),
  1103 => (x"87",x"e0",x"c3",x"02"),
  1104 => (x"1e",x"ff",x"f7",x"c0"),
  1105 => (x"c7",x"02",x"66",x"c8"),
  1106 => (x"48",x"a6",x"cc",x"87"),
  1107 => (x"87",x"c5",x"78",x"c0"),
  1108 => (x"c1",x"48",x"a6",x"cc"),
  1109 => (x"49",x"66",x"cc",x"78"),
  1110 => (x"c4",x"87",x"c2",x"e6"),
  1111 => (x"6e",x"7e",x"70",x"86"),
  1112 => (x"87",x"e9",x"c2",x"02"),
  1113 => (x"81",x"cb",x"49",x"6e"),
  1114 => (x"d0",x"49",x"69",x"97"),
  1115 => (x"d6",x"c1",x"02",x"99"),
  1116 => (x"ef",x"c2",x"c1",x"87"),
  1117 => (x"cb",x"49",x"74",x"4a"),
  1118 => (x"ce",x"e3",x"c1",x"91"),
  1119 => (x"c8",x"79",x"72",x"81"),
  1120 => (x"51",x"ff",x"c3",x"81"),
  1121 => (x"91",x"de",x"49",x"74"),
  1122 => (x"4d",x"c0",x"ed",x"c2"),
  1123 => (x"c1",x"c2",x"85",x"71"),
  1124 => (x"a5",x"c1",x"7d",x"97"),
  1125 => (x"51",x"e0",x"c0",x"49"),
  1126 => (x"97",x"f2",x"e7",x"c2"),
  1127 => (x"87",x"d2",x"02",x"bf"),
  1128 => (x"a5",x"c2",x"84",x"c1"),
  1129 => (x"f2",x"e7",x"c2",x"4b"),
  1130 => (x"fe",x"49",x"db",x"4a"),
  1131 => (x"c1",x"87",x"f9",x"fb"),
  1132 => (x"a5",x"cd",x"87",x"db"),
  1133 => (x"c1",x"51",x"c0",x"49"),
  1134 => (x"4b",x"a5",x"c2",x"84"),
  1135 => (x"49",x"cb",x"4a",x"6e"),
  1136 => (x"87",x"e4",x"fb",x"fe"),
  1137 => (x"c1",x"87",x"c6",x"c1"),
  1138 => (x"74",x"4a",x"ec",x"c0"),
  1139 => (x"c1",x"91",x"cb",x"49"),
  1140 => (x"72",x"81",x"ce",x"e3"),
  1141 => (x"f2",x"e7",x"c2",x"79"),
  1142 => (x"d8",x"02",x"bf",x"97"),
  1143 => (x"de",x"49",x"74",x"87"),
  1144 => (x"c2",x"84",x"c1",x"91"),
  1145 => (x"71",x"4b",x"c0",x"ed"),
  1146 => (x"f2",x"e7",x"c2",x"83"),
  1147 => (x"fe",x"49",x"dd",x"4a"),
  1148 => (x"d8",x"87",x"f5",x"fa"),
  1149 => (x"de",x"4b",x"74",x"87"),
  1150 => (x"c0",x"ed",x"c2",x"93"),
  1151 => (x"49",x"a3",x"cb",x"83"),
  1152 => (x"84",x"c1",x"51",x"c0"),
  1153 => (x"cb",x"4a",x"6e",x"73"),
  1154 => (x"db",x"fa",x"fe",x"49"),
  1155 => (x"48",x"66",x"c4",x"87"),
  1156 => (x"a6",x"c8",x"80",x"c1"),
  1157 => (x"03",x"ac",x"c7",x"58"),
  1158 => (x"6e",x"87",x"c5",x"c0"),
  1159 => (x"87",x"e0",x"fc",x"05"),
  1160 => (x"8e",x"f4",x"48",x"74"),
  1161 => (x"1e",x"87",x"fe",x"f5"),
  1162 => (x"4b",x"71",x"1e",x"73"),
  1163 => (x"c1",x"91",x"cb",x"49"),
  1164 => (x"c8",x"81",x"ce",x"e3"),
  1165 => (x"e2",x"c1",x"4a",x"a1"),
  1166 => (x"50",x"12",x"48",x"fe"),
  1167 => (x"c0",x"4a",x"a1",x"c9"),
  1168 => (x"12",x"48",x"ec",x"fa"),
  1169 => (x"c1",x"81",x"ca",x"50"),
  1170 => (x"11",x"48",x"ff",x"e2"),
  1171 => (x"ff",x"e2",x"c1",x"50"),
  1172 => (x"1e",x"49",x"bf",x"97"),
  1173 => (x"d3",x"f6",x"49",x"c0"),
  1174 => (x"d4",x"ec",x"c2",x"87"),
  1175 => (x"c1",x"78",x"de",x"48"),
  1176 => (x"87",x"fb",x"d5",x"49"),
  1177 => (x"87",x"c1",x"f5",x"26"),
  1178 => (x"49",x"4a",x"71",x"1e"),
  1179 => (x"e3",x"c1",x"91",x"cb"),
  1180 => (x"81",x"c8",x"81",x"ce"),
  1181 => (x"ec",x"c2",x"48",x"11"),
  1182 => (x"ec",x"c2",x"58",x"d8"),
  1183 => (x"78",x"c0",x"48",x"ec"),
  1184 => (x"da",x"d5",x"49",x"c1"),
  1185 => (x"1e",x"4f",x"26",x"87"),
  1186 => (x"fe",x"c0",x"49",x"c0"),
  1187 => (x"4f",x"26",x"87",x"ce"),
  1188 => (x"02",x"99",x"71",x"1e"),
  1189 => (x"e4",x"c1",x"87",x"d2"),
  1190 => (x"50",x"c0",x"48",x"e3"),
  1191 => (x"c9",x"c1",x"80",x"f7"),
  1192 => (x"e3",x"c1",x"40",x"e8"),
  1193 => (x"87",x"ce",x"78",x"c7"),
  1194 => (x"48",x"df",x"e4",x"c1"),
  1195 => (x"78",x"c0",x"e3",x"c1"),
  1196 => (x"ca",x"c1",x"80",x"fc"),
  1197 => (x"4f",x"26",x"78",x"c7"),
  1198 => (x"5c",x"5b",x"5e",x"0e"),
  1199 => (x"4a",x"4c",x"71",x"0e"),
  1200 => (x"e3",x"c1",x"92",x"cb"),
  1201 => (x"a2",x"c8",x"82",x"ce"),
  1202 => (x"4b",x"a2",x"c9",x"49"),
  1203 => (x"1e",x"4b",x"6b",x"97"),
  1204 => (x"1e",x"49",x"69",x"97"),
  1205 => (x"49",x"12",x"82",x"ca"),
  1206 => (x"87",x"c7",x"e7",x"c0"),
  1207 => (x"fe",x"d3",x"49",x"c0"),
  1208 => (x"c0",x"49",x"74",x"87"),
  1209 => (x"f8",x"87",x"d0",x"fb"),
  1210 => (x"87",x"fb",x"f2",x"8e"),
  1211 => (x"71",x"1e",x"73",x"1e"),
  1212 => (x"c3",x"ff",x"49",x"4b"),
  1213 => (x"fe",x"49",x"73",x"87"),
  1214 => (x"ec",x"f2",x"87",x"fe"),
  1215 => (x"1e",x"73",x"1e",x"87"),
  1216 => (x"a3",x"c6",x"4b",x"71"),
  1217 => (x"87",x"db",x"02",x"4a"),
  1218 => (x"d6",x"02",x"8a",x"c1"),
  1219 => (x"c1",x"02",x"8a",x"87"),
  1220 => (x"02",x"8a",x"87",x"da"),
  1221 => (x"8a",x"87",x"fc",x"c0"),
  1222 => (x"87",x"e1",x"c0",x"02"),
  1223 => (x"87",x"cb",x"02",x"8a"),
  1224 => (x"c7",x"87",x"db",x"c1"),
  1225 => (x"87",x"c0",x"fd",x"49"),
  1226 => (x"c2",x"87",x"de",x"c1"),
  1227 => (x"02",x"bf",x"ec",x"ec"),
  1228 => (x"48",x"87",x"cb",x"c1"),
  1229 => (x"ec",x"c2",x"88",x"c1"),
  1230 => (x"c1",x"c1",x"58",x"f0"),
  1231 => (x"f0",x"ec",x"c2",x"87"),
  1232 => (x"f9",x"c0",x"02",x"bf"),
  1233 => (x"ec",x"ec",x"c2",x"87"),
  1234 => (x"80",x"c1",x"48",x"bf"),
  1235 => (x"58",x"f0",x"ec",x"c2"),
  1236 => (x"c2",x"87",x"eb",x"c0"),
  1237 => (x"49",x"bf",x"ec",x"ec"),
  1238 => (x"ec",x"c2",x"89",x"c6"),
  1239 => (x"b7",x"c0",x"59",x"f0"),
  1240 => (x"87",x"da",x"03",x"a9"),
  1241 => (x"48",x"ec",x"ec",x"c2"),
  1242 => (x"87",x"d2",x"78",x"c0"),
  1243 => (x"bf",x"f0",x"ec",x"c2"),
  1244 => (x"c2",x"87",x"cb",x"02"),
  1245 => (x"48",x"bf",x"ec",x"ec"),
  1246 => (x"ec",x"c2",x"80",x"c6"),
  1247 => (x"49",x"c0",x"58",x"f0"),
  1248 => (x"73",x"87",x"dc",x"d1"),
  1249 => (x"ee",x"f8",x"c0",x"49"),
  1250 => (x"87",x"dd",x"f0",x"87"),
  1251 => (x"5c",x"5b",x"5e",x"0e"),
  1252 => (x"cc",x"4c",x"71",x"0e"),
  1253 => (x"4b",x"74",x"1e",x"66"),
  1254 => (x"e3",x"c1",x"93",x"cb"),
  1255 => (x"a3",x"c4",x"83",x"ce"),
  1256 => (x"fe",x"49",x"6a",x"4a"),
  1257 => (x"c1",x"87",x"d1",x"f4"),
  1258 => (x"c8",x"7b",x"e7",x"c8"),
  1259 => (x"66",x"d4",x"49",x"a3"),
  1260 => (x"49",x"a3",x"c9",x"51"),
  1261 => (x"ca",x"51",x"66",x"d8"),
  1262 => (x"66",x"dc",x"49",x"a3"),
  1263 => (x"e6",x"ef",x"26",x"51"),
  1264 => (x"5b",x"5e",x"0e",x"87"),
  1265 => (x"ff",x"0e",x"5d",x"5c"),
  1266 => (x"a6",x"d8",x"86",x"d0"),
  1267 => (x"48",x"a6",x"c4",x"59"),
  1268 => (x"80",x"c4",x"78",x"c0"),
  1269 => (x"78",x"66",x"c4",x"c1"),
  1270 => (x"78",x"c1",x"80",x"c4"),
  1271 => (x"78",x"c1",x"80",x"c4"),
  1272 => (x"48",x"f0",x"ec",x"c2"),
  1273 => (x"ec",x"c2",x"78",x"c1"),
  1274 => (x"de",x"48",x"bf",x"d4"),
  1275 => (x"87",x"cb",x"05",x"a8"),
  1276 => (x"70",x"87",x"e6",x"f3"),
  1277 => (x"59",x"a6",x"c8",x"49"),
  1278 => (x"e3",x"87",x"ec",x"ce"),
  1279 => (x"c5",x"e4",x"87",x"e3"),
  1280 => (x"87",x"d2",x"e3",x"87"),
  1281 => (x"fb",x"c0",x"4c",x"70"),
  1282 => (x"d0",x"c1",x"02",x"ac"),
  1283 => (x"05",x"66",x"d4",x"87"),
  1284 => (x"c0",x"87",x"c2",x"c1"),
  1285 => (x"1e",x"c1",x"1e",x"1e"),
  1286 => (x"1e",x"c1",x"e5",x"c1"),
  1287 => (x"eb",x"fd",x"49",x"c0"),
  1288 => (x"66",x"d0",x"c1",x"87"),
  1289 => (x"6a",x"82",x"c4",x"4a"),
  1290 => (x"74",x"81",x"c7",x"49"),
  1291 => (x"d8",x"1e",x"c1",x"51"),
  1292 => (x"c8",x"49",x"6a",x"1e"),
  1293 => (x"87",x"e2",x"e3",x"81"),
  1294 => (x"c4",x"c1",x"86",x"d8"),
  1295 => (x"a8",x"c0",x"48",x"66"),
  1296 => (x"c4",x"87",x"c7",x"01"),
  1297 => (x"78",x"c1",x"48",x"a6"),
  1298 => (x"c4",x"c1",x"87",x"ce"),
  1299 => (x"88",x"c1",x"48",x"66"),
  1300 => (x"c3",x"58",x"a6",x"cc"),
  1301 => (x"87",x"ee",x"e2",x"87"),
  1302 => (x"c2",x"48",x"a6",x"cc"),
  1303 => (x"02",x"9c",x"74",x"78"),
  1304 => (x"c4",x"87",x"c0",x"cd"),
  1305 => (x"c8",x"c1",x"48",x"66"),
  1306 => (x"cc",x"03",x"a8",x"66"),
  1307 => (x"a6",x"d8",x"87",x"f5"),
  1308 => (x"c4",x"78",x"c0",x"48"),
  1309 => (x"e1",x"78",x"c0",x"80"),
  1310 => (x"4c",x"70",x"87",x"dc"),
  1311 => (x"05",x"ac",x"d0",x"c1"),
  1312 => (x"dc",x"87",x"d8",x"c2"),
  1313 => (x"c0",x"e4",x"7e",x"66"),
  1314 => (x"c0",x"49",x"70",x"87"),
  1315 => (x"e1",x"59",x"a6",x"e0"),
  1316 => (x"4c",x"70",x"87",x"c4"),
  1317 => (x"05",x"ac",x"ec",x"c0"),
  1318 => (x"c4",x"87",x"eb",x"c1"),
  1319 => (x"91",x"cb",x"49",x"66"),
  1320 => (x"81",x"66",x"c0",x"c1"),
  1321 => (x"6a",x"4a",x"a1",x"c4"),
  1322 => (x"4a",x"a1",x"c8",x"4d"),
  1323 => (x"c1",x"52",x"66",x"dc"),
  1324 => (x"e0",x"79",x"e8",x"c9"),
  1325 => (x"4c",x"70",x"87",x"e0"),
  1326 => (x"87",x"d8",x"02",x"9c"),
  1327 => (x"02",x"ac",x"fb",x"c0"),
  1328 => (x"55",x"74",x"87",x"d2"),
  1329 => (x"70",x"87",x"cf",x"e0"),
  1330 => (x"c7",x"02",x"9c",x"4c"),
  1331 => (x"ac",x"fb",x"c0",x"87"),
  1332 => (x"87",x"ee",x"ff",x"05"),
  1333 => (x"c2",x"55",x"e0",x"c0"),
  1334 => (x"97",x"c0",x"55",x"c1"),
  1335 => (x"49",x"66",x"d4",x"7d"),
  1336 => (x"db",x"05",x"a9",x"6e"),
  1337 => (x"48",x"66",x"c4",x"87"),
  1338 => (x"04",x"a8",x"66",x"c8"),
  1339 => (x"66",x"c4",x"87",x"ca"),
  1340 => (x"c8",x"80",x"c1",x"48"),
  1341 => (x"87",x"c8",x"58",x"a6"),
  1342 => (x"c1",x"48",x"66",x"c8"),
  1343 => (x"58",x"a6",x"cc",x"88"),
  1344 => (x"87",x"d2",x"df",x"ff"),
  1345 => (x"d0",x"c1",x"4c",x"70"),
  1346 => (x"87",x"c8",x"05",x"ac"),
  1347 => (x"c1",x"48",x"66",x"d0"),
  1348 => (x"58",x"a6",x"d4",x"80"),
  1349 => (x"02",x"ac",x"d0",x"c1"),
  1350 => (x"c0",x"87",x"e8",x"fd"),
  1351 => (x"d4",x"48",x"a6",x"e0"),
  1352 => (x"66",x"dc",x"78",x"66"),
  1353 => (x"66",x"e0",x"c0",x"48"),
  1354 => (x"c8",x"c9",x"05",x"a8"),
  1355 => (x"a6",x"e4",x"c0",x"87"),
  1356 => (x"7e",x"78",x"c0",x"48"),
  1357 => (x"fb",x"c0",x"48",x"74"),
  1358 => (x"a6",x"ec",x"c0",x"88"),
  1359 => (x"02",x"98",x"70",x"58"),
  1360 => (x"48",x"87",x"cd",x"c8"),
  1361 => (x"ec",x"c0",x"88",x"cb"),
  1362 => (x"98",x"70",x"58",x"a6"),
  1363 => (x"87",x"d2",x"c1",x"02"),
  1364 => (x"c0",x"88",x"c9",x"48"),
  1365 => (x"70",x"58",x"a6",x"ec"),
  1366 => (x"db",x"c3",x"02",x"98"),
  1367 => (x"88",x"c4",x"48",x"87"),
  1368 => (x"58",x"a6",x"ec",x"c0"),
  1369 => (x"d0",x"02",x"98",x"70"),
  1370 => (x"88",x"c1",x"48",x"87"),
  1371 => (x"58",x"a6",x"ec",x"c0"),
  1372 => (x"c3",x"02",x"98",x"70"),
  1373 => (x"d1",x"c7",x"87",x"c2"),
  1374 => (x"48",x"a6",x"d8",x"87"),
  1375 => (x"ff",x"78",x"f0",x"c0"),
  1376 => (x"70",x"87",x"d3",x"dd"),
  1377 => (x"ac",x"ec",x"c0",x"4c"),
  1378 => (x"87",x"c3",x"c0",x"02"),
  1379 => (x"c0",x"5c",x"a6",x"dc"),
  1380 => (x"cd",x"02",x"ac",x"ec"),
  1381 => (x"fd",x"dc",x"ff",x"87"),
  1382 => (x"c0",x"4c",x"70",x"87"),
  1383 => (x"ff",x"05",x"ac",x"ec"),
  1384 => (x"ec",x"c0",x"87",x"f3"),
  1385 => (x"c4",x"c0",x"02",x"ac"),
  1386 => (x"e9",x"dc",x"ff",x"87"),
  1387 => (x"1e",x"66",x"d8",x"87"),
  1388 => (x"1e",x"49",x"66",x"d4"),
  1389 => (x"1e",x"49",x"66",x"d4"),
  1390 => (x"1e",x"c1",x"e5",x"c1"),
  1391 => (x"f7",x"49",x"66",x"d4"),
  1392 => (x"1e",x"c0",x"87",x"ca"),
  1393 => (x"66",x"dc",x"1e",x"ca"),
  1394 => (x"c1",x"91",x"cb",x"49"),
  1395 => (x"d8",x"81",x"66",x"d8"),
  1396 => (x"a1",x"c4",x"48",x"a6"),
  1397 => (x"bf",x"66",x"d8",x"78"),
  1398 => (x"fd",x"dc",x"ff",x"49"),
  1399 => (x"c0",x"86",x"d8",x"87"),
  1400 => (x"c1",x"06",x"a8",x"b7"),
  1401 => (x"1e",x"c1",x"87",x"c5"),
  1402 => (x"66",x"c8",x"1e",x"de"),
  1403 => (x"dc",x"ff",x"49",x"bf"),
  1404 => (x"86",x"c8",x"87",x"e8"),
  1405 => (x"c0",x"48",x"49",x"70"),
  1406 => (x"a6",x"dc",x"88",x"08"),
  1407 => (x"a8",x"b7",x"c0",x"58"),
  1408 => (x"87",x"e7",x"c0",x"06"),
  1409 => (x"dd",x"48",x"66",x"d8"),
  1410 => (x"de",x"03",x"a8",x"b7"),
  1411 => (x"49",x"bf",x"6e",x"87"),
  1412 => (x"c0",x"81",x"66",x"d8"),
  1413 => (x"66",x"d8",x"51",x"e0"),
  1414 => (x"6e",x"81",x"c1",x"49"),
  1415 => (x"c1",x"c2",x"81",x"bf"),
  1416 => (x"49",x"66",x"d8",x"51"),
  1417 => (x"bf",x"6e",x"81",x"c2"),
  1418 => (x"cc",x"51",x"c0",x"81"),
  1419 => (x"80",x"c1",x"48",x"66"),
  1420 => (x"c1",x"58",x"a6",x"d0"),
  1421 => (x"87",x"d8",x"c4",x"7e"),
  1422 => (x"87",x"cd",x"dd",x"ff"),
  1423 => (x"ff",x"58",x"a6",x"dc"),
  1424 => (x"c0",x"87",x"c6",x"dd"),
  1425 => (x"c0",x"58",x"a6",x"ec"),
  1426 => (x"c0",x"05",x"a8",x"ec"),
  1427 => (x"e8",x"c0",x"87",x"ca"),
  1428 => (x"66",x"d8",x"48",x"a6"),
  1429 => (x"87",x"c4",x"c0",x"78"),
  1430 => (x"87",x"fa",x"d9",x"ff"),
  1431 => (x"cb",x"49",x"66",x"c4"),
  1432 => (x"66",x"c0",x"c1",x"91"),
  1433 => (x"70",x"80",x"71",x"48"),
  1434 => (x"c8",x"49",x"6e",x"7e"),
  1435 => (x"ca",x"4a",x"6e",x"81"),
  1436 => (x"52",x"66",x"d8",x"82"),
  1437 => (x"4a",x"66",x"e8",x"c0"),
  1438 => (x"66",x"d8",x"82",x"c1"),
  1439 => (x"72",x"48",x"c1",x"8a"),
  1440 => (x"c1",x"4a",x"70",x"30"),
  1441 => (x"79",x"97",x"72",x"8a"),
  1442 => (x"1e",x"49",x"69",x"97"),
  1443 => (x"d7",x"49",x"66",x"dc"),
  1444 => (x"86",x"c4",x"87",x"d3"),
  1445 => (x"58",x"a6",x"f0",x"c0"),
  1446 => (x"81",x"c4",x"49",x"6e"),
  1447 => (x"e0",x"c0",x"4d",x"69"),
  1448 => (x"66",x"dc",x"48",x"66"),
  1449 => (x"c8",x"c0",x"02",x"a8"),
  1450 => (x"48",x"a6",x"d8",x"87"),
  1451 => (x"c5",x"c0",x"78",x"c0"),
  1452 => (x"48",x"a6",x"d8",x"87"),
  1453 => (x"66",x"d8",x"78",x"c1"),
  1454 => (x"1e",x"e0",x"c0",x"1e"),
  1455 => (x"d9",x"ff",x"49",x"75"),
  1456 => (x"86",x"c8",x"87",x"d8"),
  1457 => (x"b7",x"c0",x"4c",x"70"),
  1458 => (x"d4",x"c1",x"06",x"ac"),
  1459 => (x"c0",x"85",x"74",x"87"),
  1460 => (x"89",x"74",x"49",x"e0"),
  1461 => (x"df",x"c1",x"4b",x"75"),
  1462 => (x"fe",x"71",x"4a",x"dc"),
  1463 => (x"c2",x"87",x"c9",x"e7"),
  1464 => (x"66",x"e4",x"c0",x"85"),
  1465 => (x"c0",x"80",x"c1",x"48"),
  1466 => (x"c0",x"58",x"a6",x"e8"),
  1467 => (x"c1",x"49",x"66",x"ec"),
  1468 => (x"02",x"a9",x"70",x"81"),
  1469 => (x"d8",x"87",x"c8",x"c0"),
  1470 => (x"78",x"c0",x"48",x"a6"),
  1471 => (x"d8",x"87",x"c5",x"c0"),
  1472 => (x"78",x"c1",x"48",x"a6"),
  1473 => (x"c2",x"1e",x"66",x"d8"),
  1474 => (x"e0",x"c0",x"49",x"a4"),
  1475 => (x"70",x"88",x"71",x"48"),
  1476 => (x"49",x"75",x"1e",x"49"),
  1477 => (x"87",x"c2",x"d8",x"ff"),
  1478 => (x"b7",x"c0",x"86",x"c8"),
  1479 => (x"c0",x"ff",x"01",x"a8"),
  1480 => (x"66",x"e4",x"c0",x"87"),
  1481 => (x"87",x"d1",x"c0",x"02"),
  1482 => (x"81",x"c9",x"49",x"6e"),
  1483 => (x"51",x"66",x"e4",x"c0"),
  1484 => (x"ca",x"c1",x"48",x"6e"),
  1485 => (x"cc",x"c0",x"78",x"f8"),
  1486 => (x"c9",x"49",x"6e",x"87"),
  1487 => (x"6e",x"51",x"c2",x"81"),
  1488 => (x"ec",x"cb",x"c1",x"48"),
  1489 => (x"c0",x"7e",x"c1",x"78"),
  1490 => (x"d6",x"ff",x"87",x"c6"),
  1491 => (x"4c",x"70",x"87",x"f8"),
  1492 => (x"f5",x"c0",x"02",x"6e"),
  1493 => (x"48",x"66",x"c4",x"87"),
  1494 => (x"04",x"a8",x"66",x"c8"),
  1495 => (x"c4",x"87",x"cb",x"c0"),
  1496 => (x"80",x"c1",x"48",x"66"),
  1497 => (x"c0",x"58",x"a6",x"c8"),
  1498 => (x"66",x"c8",x"87",x"e0"),
  1499 => (x"cc",x"88",x"c1",x"48"),
  1500 => (x"d5",x"c0",x"58",x"a6"),
  1501 => (x"ac",x"c6",x"c1",x"87"),
  1502 => (x"87",x"c8",x"c0",x"05"),
  1503 => (x"c1",x"48",x"66",x"cc"),
  1504 => (x"58",x"a6",x"d0",x"80"),
  1505 => (x"87",x"fe",x"d5",x"ff"),
  1506 => (x"66",x"d0",x"4c",x"70"),
  1507 => (x"d4",x"80",x"c1",x"48"),
  1508 => (x"9c",x"74",x"58",x"a6"),
  1509 => (x"87",x"cb",x"c0",x"02"),
  1510 => (x"c1",x"48",x"66",x"c4"),
  1511 => (x"04",x"a8",x"66",x"c8"),
  1512 => (x"ff",x"87",x"cb",x"f3"),
  1513 => (x"c4",x"87",x"d6",x"d5"),
  1514 => (x"a8",x"c7",x"48",x"66"),
  1515 => (x"87",x"e5",x"c0",x"03"),
  1516 => (x"48",x"f0",x"ec",x"c2"),
  1517 => (x"66",x"c4",x"78",x"c0"),
  1518 => (x"c1",x"91",x"cb",x"49"),
  1519 => (x"c4",x"81",x"66",x"c0"),
  1520 => (x"4a",x"6a",x"4a",x"a1"),
  1521 => (x"c4",x"79",x"52",x"c0"),
  1522 => (x"80",x"c1",x"48",x"66"),
  1523 => (x"c7",x"58",x"a6",x"c8"),
  1524 => (x"db",x"ff",x"04",x"a8"),
  1525 => (x"8e",x"d0",x"ff",x"87"),
  1526 => (x"87",x"c9",x"df",x"ff"),
  1527 => (x"1e",x"00",x"20",x"3a"),
  1528 => (x"4b",x"71",x"1e",x"73"),
  1529 => (x"87",x"c6",x"02",x"9b"),
  1530 => (x"48",x"ec",x"ec",x"c2"),
  1531 => (x"1e",x"c7",x"78",x"c0"),
  1532 => (x"bf",x"ec",x"ec",x"c2"),
  1533 => (x"e3",x"c1",x"1e",x"49"),
  1534 => (x"ec",x"c2",x"1e",x"ce"),
  1535 => (x"ee",x"49",x"bf",x"d4"),
  1536 => (x"86",x"cc",x"87",x"ff"),
  1537 => (x"bf",x"d4",x"ec",x"c2"),
  1538 => (x"87",x"c4",x"ea",x"49"),
  1539 => (x"c8",x"02",x"9b",x"73"),
  1540 => (x"ce",x"e3",x"c1",x"87"),
  1541 => (x"f0",x"e7",x"c0",x"49"),
  1542 => (x"cc",x"de",x"ff",x"87"),
  1543 => (x"e2",x"c1",x"1e",x"87"),
  1544 => (x"50",x"c0",x"48",x"fe"),
  1545 => (x"bf",x"f1",x"e4",x"c1"),
  1546 => (x"c0",x"da",x"ff",x"49"),
  1547 => (x"26",x"48",x"c0",x"87"),
  1548 => (x"eb",x"c7",x"1e",x"4f"),
  1549 => (x"fe",x"49",x"c1",x"87"),
  1550 => (x"ea",x"fe",x"87",x"e5"),
  1551 => (x"98",x"70",x"87",x"df"),
  1552 => (x"fe",x"87",x"cd",x"02"),
  1553 => (x"70",x"87",x"da",x"f3"),
  1554 => (x"87",x"c4",x"02",x"98"),
  1555 => (x"87",x"c2",x"4a",x"c1"),
  1556 => (x"9a",x"72",x"4a",x"c0"),
  1557 => (x"c0",x"87",x"ce",x"05"),
  1558 => (x"c5",x"e2",x"c1",x"1e"),
  1559 => (x"c0",x"f3",x"c0",x"49"),
  1560 => (x"fe",x"86",x"c4",x"87"),
  1561 => (x"e8",x"fc",x"c0",x"87"),
  1562 => (x"c1",x"1e",x"c0",x"87"),
  1563 => (x"c0",x"49",x"d0",x"e2"),
  1564 => (x"c0",x"87",x"ee",x"f2"),
  1565 => (x"87",x"e5",x"fe",x"1e"),
  1566 => (x"f2",x"c0",x"49",x"70"),
  1567 => (x"de",x"c3",x"87",x"e3"),
  1568 => (x"26",x"8e",x"f8",x"87"),
  1569 => (x"20",x"44",x"53",x"4f"),
  1570 => (x"6c",x"69",x"61",x"66"),
  1571 => (x"00",x"2e",x"64",x"65"),
  1572 => (x"74",x"6f",x"6f",x"42"),
  1573 => (x"2e",x"67",x"6e",x"69"),
  1574 => (x"1e",x"00",x"2e",x"2e"),
  1575 => (x"87",x"c5",x"ea",x"c0"),
  1576 => (x"87",x"f3",x"f5",x"c0"),
  1577 => (x"4f",x"26",x"87",x"f6"),
  1578 => (x"ec",x"ec",x"c2",x"1e"),
  1579 => (x"c2",x"78",x"c0",x"48"),
  1580 => (x"c0",x"48",x"d4",x"ec"),
  1581 => (x"87",x"f9",x"fd",x"78"),
  1582 => (x"48",x"c0",x"87",x"e1"),
  1583 => (x"00",x"00",x"4f",x"26"),
  1584 => (x"78",x"45",x"20",x"80"),
  1585 => (x"80",x"00",x"74",x"69"),
  1586 => (x"63",x"61",x"42",x"20"),
  1587 => (x"12",x"68",x"00",x"6b"),
  1588 => (x"2b",x"40",x"00",x"00"),
  1589 => (x"00",x"00",x"00",x"00"),
  1590 => (x"00",x"12",x"68",x"00"),
  1591 => (x"00",x"2b",x"5e",x"00"),
  1592 => (x"00",x"00",x"00",x"00"),
  1593 => (x"00",x"00",x"12",x"68"),
  1594 => (x"00",x"00",x"2b",x"7c"),
  1595 => (x"68",x"00",x"00",x"00"),
  1596 => (x"9a",x"00",x"00",x"12"),
  1597 => (x"00",x"00",x"00",x"2b"),
  1598 => (x"12",x"68",x"00",x"00"),
  1599 => (x"2b",x"b8",x"00",x"00"),
  1600 => (x"00",x"00",x"00",x"00"),
  1601 => (x"00",x"12",x"68",x"00"),
  1602 => (x"00",x"2b",x"d6",x"00"),
  1603 => (x"00",x"00",x"00",x"00"),
  1604 => (x"00",x"00",x"12",x"68"),
  1605 => (x"00",x"00",x"2b",x"f4"),
  1606 => (x"68",x"00",x"00",x"00"),
  1607 => (x"00",x"00",x"00",x"12"),
  1608 => (x"00",x"00",x"00",x"00"),
  1609 => (x"12",x"fd",x"00",x"00"),
  1610 => (x"00",x"00",x"00",x"00"),
  1611 => (x"00",x"00",x"00",x"00"),
  1612 => (x"00",x"19",x"35",x"00"),
  1613 => (x"34",x"36",x"43",x"00"),
  1614 => (x"20",x"20",x"20",x"20"),
  1615 => (x"4d",x"4f",x"52",x"20"),
  1616 => (x"61",x"6f",x"4c",x"00"),
  1617 => (x"2e",x"2a",x"20",x"64"),
  1618 => (x"f0",x"fe",x"1e",x"00"),
  1619 => (x"cd",x"78",x"c0",x"48"),
  1620 => (x"26",x"09",x"79",x"09"),
  1621 => (x"fe",x"1e",x"1e",x"4f"),
  1622 => (x"48",x"7e",x"bf",x"f0"),
  1623 => (x"1e",x"4f",x"26",x"26"),
  1624 => (x"c1",x"48",x"f0",x"fe"),
  1625 => (x"1e",x"4f",x"26",x"78"),
  1626 => (x"c0",x"48",x"f0",x"fe"),
  1627 => (x"1e",x"4f",x"26",x"78"),
  1628 => (x"52",x"c0",x"4a",x"71"),
  1629 => (x"0e",x"4f",x"26",x"52"),
  1630 => (x"5d",x"5c",x"5b",x"5e"),
  1631 => (x"71",x"86",x"f4",x"0e"),
  1632 => (x"7e",x"6d",x"97",x"4d"),
  1633 => (x"97",x"4c",x"a5",x"c1"),
  1634 => (x"a6",x"c8",x"48",x"6c"),
  1635 => (x"c4",x"48",x"6e",x"58"),
  1636 => (x"c5",x"05",x"a8",x"66"),
  1637 => (x"c0",x"48",x"ff",x"87"),
  1638 => (x"ca",x"ff",x"87",x"e6"),
  1639 => (x"49",x"a5",x"c2",x"87"),
  1640 => (x"71",x"4b",x"6c",x"97"),
  1641 => (x"6b",x"97",x"4b",x"a3"),
  1642 => (x"7e",x"6c",x"97",x"4b"),
  1643 => (x"80",x"c1",x"48",x"6e"),
  1644 => (x"c7",x"58",x"a6",x"c8"),
  1645 => (x"58",x"a6",x"cc",x"98"),
  1646 => (x"fe",x"7c",x"97",x"70"),
  1647 => (x"48",x"73",x"87",x"e1"),
  1648 => (x"4d",x"26",x"8e",x"f4"),
  1649 => (x"4b",x"26",x"4c",x"26"),
  1650 => (x"5e",x"0e",x"4f",x"26"),
  1651 => (x"f4",x"0e",x"5c",x"5b"),
  1652 => (x"d8",x"4c",x"71",x"86"),
  1653 => (x"ff",x"c3",x"4a",x"66"),
  1654 => (x"4b",x"a4",x"c2",x"9a"),
  1655 => (x"73",x"49",x"6c",x"97"),
  1656 => (x"51",x"72",x"49",x"a1"),
  1657 => (x"6e",x"7e",x"6c",x"97"),
  1658 => (x"c8",x"80",x"c1",x"48"),
  1659 => (x"98",x"c7",x"58",x"a6"),
  1660 => (x"70",x"58",x"a6",x"cc"),
  1661 => (x"ff",x"8e",x"f4",x"54"),
  1662 => (x"1e",x"1e",x"87",x"ca"),
  1663 => (x"e0",x"87",x"e8",x"fd"),
  1664 => (x"c0",x"49",x"4a",x"bf"),
  1665 => (x"02",x"99",x"c0",x"e0"),
  1666 => (x"1e",x"72",x"87",x"cb"),
  1667 => (x"49",x"d2",x"f0",x"c2"),
  1668 => (x"c4",x"87",x"f7",x"fe"),
  1669 => (x"87",x"fd",x"fc",x"86"),
  1670 => (x"c2",x"fd",x"7e",x"70"),
  1671 => (x"4f",x"26",x"26",x"87"),
  1672 => (x"d2",x"f0",x"c2",x"1e"),
  1673 => (x"87",x"c7",x"fd",x"49"),
  1674 => (x"49",x"fa",x"e7",x"c1"),
  1675 => (x"c4",x"87",x"da",x"fc"),
  1676 => (x"4f",x"26",x"87",x"c8"),
  1677 => (x"48",x"d0",x"ff",x"1e"),
  1678 => (x"ff",x"78",x"e1",x"c8"),
  1679 => (x"78",x"c5",x"48",x"d4"),
  1680 => (x"c3",x"02",x"66",x"c4"),
  1681 => (x"78",x"e0",x"c3",x"87"),
  1682 => (x"c6",x"02",x"66",x"c8"),
  1683 => (x"48",x"d4",x"ff",x"87"),
  1684 => (x"ff",x"78",x"f0",x"c3"),
  1685 => (x"78",x"71",x"48",x"d4"),
  1686 => (x"c8",x"48",x"d0",x"ff"),
  1687 => (x"e0",x"c0",x"78",x"e1"),
  1688 => (x"0e",x"4f",x"26",x"78"),
  1689 => (x"0e",x"5c",x"5b",x"5e"),
  1690 => (x"f0",x"c2",x"4c",x"71"),
  1691 => (x"c6",x"fc",x"49",x"d2"),
  1692 => (x"c0",x"4a",x"70",x"87"),
  1693 => (x"c2",x"04",x"aa",x"b7"),
  1694 => (x"e0",x"c3",x"87",x"e3"),
  1695 => (x"87",x"c9",x"05",x"aa"),
  1696 => (x"48",x"ed",x"ec",x"c1"),
  1697 => (x"d4",x"c2",x"78",x"c1"),
  1698 => (x"aa",x"f0",x"c3",x"87"),
  1699 => (x"c1",x"87",x"c9",x"05"),
  1700 => (x"c1",x"48",x"e9",x"ec"),
  1701 => (x"87",x"f5",x"c1",x"78"),
  1702 => (x"bf",x"ed",x"ec",x"c1"),
  1703 => (x"72",x"87",x"c7",x"02"),
  1704 => (x"b3",x"c0",x"c2",x"4b"),
  1705 => (x"4b",x"72",x"87",x"c2"),
  1706 => (x"d1",x"05",x"9c",x"74"),
  1707 => (x"e9",x"ec",x"c1",x"87"),
  1708 => (x"ec",x"c1",x"1e",x"bf"),
  1709 => (x"72",x"1e",x"bf",x"ed"),
  1710 => (x"87",x"f8",x"fd",x"49"),
  1711 => (x"ec",x"c1",x"86",x"c8"),
  1712 => (x"c0",x"02",x"bf",x"e9"),
  1713 => (x"49",x"73",x"87",x"e0"),
  1714 => (x"91",x"29",x"b7",x"c4"),
  1715 => (x"81",x"c9",x"ee",x"c1"),
  1716 => (x"9a",x"cf",x"4a",x"73"),
  1717 => (x"48",x"c1",x"92",x"c2"),
  1718 => (x"4a",x"70",x"30",x"72"),
  1719 => (x"48",x"72",x"ba",x"ff"),
  1720 => (x"79",x"70",x"98",x"69"),
  1721 => (x"49",x"73",x"87",x"db"),
  1722 => (x"91",x"29",x"b7",x"c4"),
  1723 => (x"81",x"c9",x"ee",x"c1"),
  1724 => (x"9a",x"cf",x"4a",x"73"),
  1725 => (x"48",x"c3",x"92",x"c2"),
  1726 => (x"4a",x"70",x"30",x"72"),
  1727 => (x"70",x"b0",x"69",x"48"),
  1728 => (x"ed",x"ec",x"c1",x"79"),
  1729 => (x"c1",x"78",x"c0",x"48"),
  1730 => (x"c0",x"48",x"e9",x"ec"),
  1731 => (x"d2",x"f0",x"c2",x"78"),
  1732 => (x"87",x"e3",x"f9",x"49"),
  1733 => (x"b7",x"c0",x"4a",x"70"),
  1734 => (x"dd",x"fd",x"03",x"aa"),
  1735 => (x"c2",x"48",x"c0",x"87"),
  1736 => (x"26",x"4d",x"26",x"87"),
  1737 => (x"26",x"4b",x"26",x"4c"),
  1738 => (x"00",x"00",x"00",x"4f"),
  1739 => (x"00",x"00",x"00",x"00"),
  1740 => (x"4a",x"71",x"1e",x"00"),
  1741 => (x"87",x"eb",x"fc",x"49"),
  1742 => (x"c0",x"1e",x"4f",x"26"),
  1743 => (x"c4",x"49",x"72",x"4a"),
  1744 => (x"c9",x"ee",x"c1",x"91"),
  1745 => (x"c1",x"79",x"c0",x"81"),
  1746 => (x"aa",x"b7",x"d0",x"82"),
  1747 => (x"26",x"87",x"ee",x"04"),
  1748 => (x"5b",x"5e",x"0e",x"4f"),
  1749 => (x"71",x"0e",x"5d",x"5c"),
  1750 => (x"87",x"cb",x"f8",x"4d"),
  1751 => (x"b7",x"c4",x"4a",x"75"),
  1752 => (x"ee",x"c1",x"92",x"2a"),
  1753 => (x"4c",x"75",x"82",x"c9"),
  1754 => (x"94",x"c2",x"9c",x"cf"),
  1755 => (x"74",x"4b",x"49",x"6a"),
  1756 => (x"c2",x"9b",x"c3",x"2b"),
  1757 => (x"70",x"30",x"74",x"48"),
  1758 => (x"74",x"bc",x"ff",x"4c"),
  1759 => (x"70",x"98",x"71",x"48"),
  1760 => (x"87",x"db",x"f7",x"7a"),
  1761 => (x"d8",x"fe",x"48",x"73"),
  1762 => (x"00",x"00",x"00",x"87"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"00",x"00",x"00"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"00",x"00",x"00",x"00"),
  1776 => (x"00",x"00",x"00",x"00"),
  1777 => (x"00",x"00",x"00",x"00"),
  1778 => (x"d0",x"ff",x"1e",x"00"),
  1779 => (x"78",x"e1",x"c8",x"48"),
  1780 => (x"d4",x"ff",x"48",x"71"),
  1781 => (x"4f",x"26",x"78",x"08"),
  1782 => (x"48",x"d0",x"ff",x"1e"),
  1783 => (x"71",x"78",x"e1",x"c8"),
  1784 => (x"08",x"d4",x"ff",x"48"),
  1785 => (x"48",x"66",x"c4",x"78"),
  1786 => (x"78",x"08",x"d4",x"ff"),
  1787 => (x"71",x"1e",x"4f",x"26"),
  1788 => (x"49",x"66",x"c4",x"4a"),
  1789 => (x"ff",x"49",x"72",x"1e"),
  1790 => (x"d0",x"ff",x"87",x"de"),
  1791 => (x"78",x"e0",x"c0",x"48"),
  1792 => (x"1e",x"4f",x"26",x"26"),
  1793 => (x"4b",x"71",x"1e",x"73"),
  1794 => (x"1e",x"49",x"66",x"c8"),
  1795 => (x"e0",x"c1",x"4a",x"73"),
  1796 => (x"d9",x"ff",x"49",x"a2"),
  1797 => (x"87",x"c4",x"26",x"87"),
  1798 => (x"4c",x"26",x"4d",x"26"),
  1799 => (x"4f",x"26",x"4b",x"26"),
  1800 => (x"4a",x"d4",x"ff",x"1e"),
  1801 => (x"ff",x"7a",x"ff",x"c3"),
  1802 => (x"e1",x"c8",x"48",x"d0"),
  1803 => (x"c2",x"7a",x"de",x"78"),
  1804 => (x"7a",x"bf",x"dc",x"f0"),
  1805 => (x"28",x"c8",x"48",x"49"),
  1806 => (x"48",x"71",x"7a",x"70"),
  1807 => (x"7a",x"70",x"28",x"d0"),
  1808 => (x"28",x"d8",x"48",x"71"),
  1809 => (x"f0",x"c2",x"7a",x"70"),
  1810 => (x"49",x"7a",x"bf",x"e0"),
  1811 => (x"70",x"28",x"c8",x"48"),
  1812 => (x"d0",x"48",x"71",x"7a"),
  1813 => (x"71",x"7a",x"70",x"28"),
  1814 => (x"70",x"28",x"d8",x"48"),
  1815 => (x"48",x"d0",x"ff",x"7a"),
  1816 => (x"26",x"78",x"e0",x"c0"),
  1817 => (x"1e",x"73",x"1e",x"4f"),
  1818 => (x"f0",x"c2",x"4a",x"71"),
  1819 => (x"72",x"4b",x"bf",x"dc"),
  1820 => (x"aa",x"e0",x"c0",x"2b"),
  1821 => (x"72",x"87",x"ce",x"04"),
  1822 => (x"89",x"e0",x"c0",x"49"),
  1823 => (x"bf",x"e0",x"f0",x"c2"),
  1824 => (x"cf",x"2b",x"71",x"4b"),
  1825 => (x"49",x"e0",x"c0",x"87"),
  1826 => (x"f0",x"c2",x"89",x"72"),
  1827 => (x"71",x"48",x"bf",x"e0"),
  1828 => (x"b3",x"49",x"70",x"30"),
  1829 => (x"73",x"9b",x"66",x"c8"),
  1830 => (x"26",x"87",x"c4",x"48"),
  1831 => (x"26",x"4c",x"26",x"4d"),
  1832 => (x"0e",x"4f",x"26",x"4b"),
  1833 => (x"5d",x"5c",x"5b",x"5e"),
  1834 => (x"71",x"86",x"ec",x"0e"),
  1835 => (x"dc",x"f0",x"c2",x"4b"),
  1836 => (x"73",x"4c",x"7e",x"bf"),
  1837 => (x"ab",x"e0",x"c0",x"2c"),
  1838 => (x"87",x"e0",x"c0",x"04"),
  1839 => (x"c0",x"48",x"a6",x"c4"),
  1840 => (x"c0",x"49",x"73",x"78"),
  1841 => (x"4a",x"71",x"89",x"e0"),
  1842 => (x"48",x"66",x"e4",x"c0"),
  1843 => (x"a6",x"cc",x"30",x"72"),
  1844 => (x"e0",x"f0",x"c2",x"58"),
  1845 => (x"71",x"4c",x"4d",x"bf"),
  1846 => (x"87",x"e4",x"c0",x"2c"),
  1847 => (x"e4",x"c0",x"49",x"73"),
  1848 => (x"30",x"71",x"48",x"66"),
  1849 => (x"c0",x"58",x"a6",x"c8"),
  1850 => (x"89",x"73",x"49",x"e0"),
  1851 => (x"48",x"66",x"e4",x"c0"),
  1852 => (x"a6",x"cc",x"28",x"71"),
  1853 => (x"e0",x"f0",x"c2",x"58"),
  1854 => (x"71",x"48",x"4d",x"bf"),
  1855 => (x"b4",x"49",x"70",x"30"),
  1856 => (x"9c",x"66",x"e4",x"c0"),
  1857 => (x"e8",x"c0",x"84",x"c1"),
  1858 => (x"c2",x"04",x"ac",x"66"),
  1859 => (x"c0",x"4c",x"c0",x"87"),
  1860 => (x"d3",x"04",x"ab",x"e0"),
  1861 => (x"48",x"a6",x"cc",x"87"),
  1862 => (x"49",x"73",x"78",x"c0"),
  1863 => (x"74",x"89",x"e0",x"c0"),
  1864 => (x"d4",x"30",x"71",x"48"),
  1865 => (x"87",x"d5",x"58",x"a6"),
  1866 => (x"48",x"74",x"49",x"73"),
  1867 => (x"a6",x"d0",x"30",x"71"),
  1868 => (x"49",x"e0",x"c0",x"58"),
  1869 => (x"48",x"74",x"89",x"73"),
  1870 => (x"a6",x"d4",x"28",x"71"),
  1871 => (x"4a",x"66",x"c4",x"58"),
  1872 => (x"9a",x"6e",x"ba",x"ff"),
  1873 => (x"ff",x"49",x"66",x"c8"),
  1874 => (x"72",x"99",x"75",x"b9"),
  1875 => (x"b0",x"66",x"cc",x"48"),
  1876 => (x"58",x"e0",x"f0",x"c2"),
  1877 => (x"66",x"d0",x"48",x"71"),
  1878 => (x"e4",x"f0",x"c2",x"b0"),
  1879 => (x"87",x"c0",x"fb",x"58"),
  1880 => (x"f6",x"fc",x"8e",x"ec"),
  1881 => (x"d0",x"ff",x"1e",x"87"),
  1882 => (x"78",x"c9",x"c8",x"48"),
  1883 => (x"d4",x"ff",x"48",x"71"),
  1884 => (x"4f",x"26",x"78",x"08"),
  1885 => (x"49",x"4a",x"71",x"1e"),
  1886 => (x"d0",x"ff",x"87",x"eb"),
  1887 => (x"26",x"78",x"c8",x"48"),
  1888 => (x"1e",x"73",x"1e",x"4f"),
  1889 => (x"f0",x"c2",x"4b",x"71"),
  1890 => (x"c3",x"02",x"bf",x"f0"),
  1891 => (x"87",x"eb",x"c2",x"87"),
  1892 => (x"c8",x"48",x"d0",x"ff"),
  1893 => (x"49",x"73",x"78",x"c9"),
  1894 => (x"ff",x"b1",x"e0",x"c0"),
  1895 => (x"78",x"71",x"48",x"d4"),
  1896 => (x"48",x"e4",x"f0",x"c2"),
  1897 => (x"66",x"c8",x"78",x"c0"),
  1898 => (x"c3",x"87",x"c5",x"02"),
  1899 => (x"87",x"c2",x"49",x"ff"),
  1900 => (x"f0",x"c2",x"49",x"c0"),
  1901 => (x"66",x"cc",x"59",x"ec"),
  1902 => (x"c5",x"87",x"c6",x"02"),
  1903 => (x"c4",x"4a",x"d5",x"d5"),
  1904 => (x"ff",x"ff",x"cf",x"87"),
  1905 => (x"f0",x"f0",x"c2",x"4a"),
  1906 => (x"f0",x"f0",x"c2",x"5a"),
  1907 => (x"c4",x"78",x"c1",x"48"),
  1908 => (x"26",x"4d",x"26",x"87"),
  1909 => (x"26",x"4b",x"26",x"4c"),
  1910 => (x"5b",x"5e",x"0e",x"4f"),
  1911 => (x"71",x"0e",x"5d",x"5c"),
  1912 => (x"ec",x"f0",x"c2",x"4a"),
  1913 => (x"9a",x"72",x"4c",x"bf"),
  1914 => (x"49",x"87",x"cb",x"02"),
  1915 => (x"f5",x"c1",x"91",x"c8"),
  1916 => (x"83",x"71",x"4b",x"f7"),
  1917 => (x"f9",x"c1",x"87",x"c4"),
  1918 => (x"4d",x"c0",x"4b",x"f7"),
  1919 => (x"99",x"74",x"49",x"13"),
  1920 => (x"bf",x"e8",x"f0",x"c2"),
  1921 => (x"48",x"d4",x"ff",x"b9"),
  1922 => (x"b7",x"c1",x"78",x"71"),
  1923 => (x"b7",x"c8",x"85",x"2c"),
  1924 => (x"87",x"e8",x"04",x"ad"),
  1925 => (x"bf",x"e4",x"f0",x"c2"),
  1926 => (x"c2",x"80",x"c8",x"48"),
  1927 => (x"fe",x"58",x"e8",x"f0"),
  1928 => (x"73",x"1e",x"87",x"ef"),
  1929 => (x"13",x"4b",x"71",x"1e"),
  1930 => (x"cb",x"02",x"9a",x"4a"),
  1931 => (x"fe",x"49",x"72",x"87"),
  1932 => (x"4a",x"13",x"87",x"e7"),
  1933 => (x"87",x"f5",x"05",x"9a"),
  1934 => (x"1e",x"87",x"da",x"fe"),
  1935 => (x"bf",x"e4",x"f0",x"c2"),
  1936 => (x"e4",x"f0",x"c2",x"49"),
  1937 => (x"78",x"a1",x"c1",x"48"),
  1938 => (x"a9",x"b7",x"c0",x"c4"),
  1939 => (x"ff",x"87",x"db",x"03"),
  1940 => (x"f0",x"c2",x"48",x"d4"),
  1941 => (x"c2",x"78",x"bf",x"e8"),
  1942 => (x"49",x"bf",x"e4",x"f0"),
  1943 => (x"48",x"e4",x"f0",x"c2"),
  1944 => (x"c4",x"78",x"a1",x"c1"),
  1945 => (x"04",x"a9",x"b7",x"c0"),
  1946 => (x"d0",x"ff",x"87",x"e5"),
  1947 => (x"c2",x"78",x"c8",x"48"),
  1948 => (x"c0",x"48",x"f0",x"f0"),
  1949 => (x"00",x"4f",x"26",x"78"),
  1950 => (x"00",x"00",x"00",x"00"),
  1951 => (x"00",x"00",x"00",x"00"),
  1952 => (x"5f",x"5f",x"00",x"00"),
  1953 => (x"00",x"00",x"00",x"00"),
  1954 => (x"03",x"00",x"03",x"03"),
  1955 => (x"14",x"00",x"00",x"03"),
  1956 => (x"7f",x"14",x"7f",x"7f"),
  1957 => (x"00",x"00",x"14",x"7f"),
  1958 => (x"6b",x"6b",x"2e",x"24"),
  1959 => (x"4c",x"00",x"12",x"3a"),
  1960 => (x"6c",x"18",x"36",x"6a"),
  1961 => (x"30",x"00",x"32",x"56"),
  1962 => (x"77",x"59",x"4f",x"7e"),
  1963 => (x"00",x"40",x"68",x"3a"),
  1964 => (x"03",x"07",x"04",x"00"),
  1965 => (x"00",x"00",x"00",x"00"),
  1966 => (x"63",x"3e",x"1c",x"00"),
  1967 => (x"00",x"00",x"00",x"41"),
  1968 => (x"3e",x"63",x"41",x"00"),
  1969 => (x"08",x"00",x"00",x"1c"),
  1970 => (x"1c",x"1c",x"3e",x"2a"),
  1971 => (x"00",x"08",x"2a",x"3e"),
  1972 => (x"3e",x"3e",x"08",x"08"),
  1973 => (x"00",x"00",x"08",x"08"),
  1974 => (x"60",x"e0",x"80",x"00"),
  1975 => (x"00",x"00",x"00",x"00"),
  1976 => (x"08",x"08",x"08",x"08"),
  1977 => (x"00",x"00",x"08",x"08"),
  1978 => (x"60",x"60",x"00",x"00"),
  1979 => (x"40",x"00",x"00",x"00"),
  1980 => (x"0c",x"18",x"30",x"60"),
  1981 => (x"00",x"01",x"03",x"06"),
  1982 => (x"4d",x"59",x"7f",x"3e"),
  1983 => (x"00",x"00",x"3e",x"7f"),
  1984 => (x"7f",x"7f",x"06",x"04"),
  1985 => (x"00",x"00",x"00",x"00"),
  1986 => (x"59",x"71",x"63",x"42"),
  1987 => (x"00",x"00",x"46",x"4f"),
  1988 => (x"49",x"49",x"63",x"22"),
  1989 => (x"18",x"00",x"36",x"7f"),
  1990 => (x"7f",x"13",x"16",x"1c"),
  1991 => (x"00",x"00",x"10",x"7f"),
  1992 => (x"45",x"45",x"67",x"27"),
  1993 => (x"00",x"00",x"39",x"7d"),
  1994 => (x"49",x"4b",x"7e",x"3c"),
  1995 => (x"00",x"00",x"30",x"79"),
  1996 => (x"79",x"71",x"01",x"01"),
  1997 => (x"00",x"00",x"07",x"0f"),
  1998 => (x"49",x"49",x"7f",x"36"),
  1999 => (x"00",x"00",x"36",x"7f"),
  2000 => (x"69",x"49",x"4f",x"06"),
  2001 => (x"00",x"00",x"1e",x"3f"),
  2002 => (x"66",x"66",x"00",x"00"),
  2003 => (x"00",x"00",x"00",x"00"),
  2004 => (x"66",x"e6",x"80",x"00"),
  2005 => (x"00",x"00",x"00",x"00"),
  2006 => (x"14",x"14",x"08",x"08"),
  2007 => (x"00",x"00",x"22",x"22"),
  2008 => (x"14",x"14",x"14",x"14"),
  2009 => (x"00",x"00",x"14",x"14"),
  2010 => (x"14",x"14",x"22",x"22"),
  2011 => (x"00",x"00",x"08",x"08"),
  2012 => (x"59",x"51",x"03",x"02"),
  2013 => (x"3e",x"00",x"06",x"0f"),
  2014 => (x"55",x"5d",x"41",x"7f"),
  2015 => (x"00",x"00",x"1e",x"1f"),
  2016 => (x"09",x"09",x"7f",x"7e"),
  2017 => (x"00",x"00",x"7e",x"7f"),
  2018 => (x"49",x"49",x"7f",x"7f"),
  2019 => (x"00",x"00",x"36",x"7f"),
  2020 => (x"41",x"63",x"3e",x"1c"),
  2021 => (x"00",x"00",x"41",x"41"),
  2022 => (x"63",x"41",x"7f",x"7f"),
  2023 => (x"00",x"00",x"1c",x"3e"),
  2024 => (x"49",x"49",x"7f",x"7f"),
  2025 => (x"00",x"00",x"41",x"41"),
  2026 => (x"09",x"09",x"7f",x"7f"),
  2027 => (x"00",x"00",x"01",x"01"),
  2028 => (x"49",x"41",x"7f",x"3e"),
  2029 => (x"00",x"00",x"7a",x"7b"),
  2030 => (x"08",x"08",x"7f",x"7f"),
  2031 => (x"00",x"00",x"7f",x"7f"),
  2032 => (x"7f",x"7f",x"41",x"00"),
  2033 => (x"00",x"00",x"00",x"41"),
  2034 => (x"40",x"40",x"60",x"20"),
  2035 => (x"7f",x"00",x"3f",x"7f"),
  2036 => (x"36",x"1c",x"08",x"7f"),
  2037 => (x"00",x"00",x"41",x"63"),
  2038 => (x"40",x"40",x"7f",x"7f"),
  2039 => (x"7f",x"00",x"40",x"40"),
  2040 => (x"06",x"0c",x"06",x"7f"),
  2041 => (x"7f",x"00",x"7f",x"7f"),
  2042 => (x"18",x"0c",x"06",x"7f"),
  2043 => (x"00",x"00",x"7f",x"7f"),
  2044 => (x"41",x"41",x"7f",x"3e"),
  2045 => (x"00",x"00",x"3e",x"7f"),
  2046 => (x"09",x"09",x"7f",x"7f"),
  2047 => (x"3e",x"00",x"06",x"0f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

