
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"00",x"40",x"7e"),
     1 => (x"19",x"09",x"7f",x"7f"),
     2 => (x"00",x"00",x"66",x"7f"),
     3 => (x"59",x"4d",x"6f",x"26"),
     4 => (x"00",x"00",x"32",x"7b"),
     5 => (x"7f",x"7f",x"01",x"01"),
     6 => (x"00",x"00",x"01",x"01"),
     7 => (x"40",x"40",x"7f",x"3f"),
     8 => (x"00",x"00",x"3f",x"7f"),
     9 => (x"70",x"70",x"3f",x"0f"),
    10 => (x"7f",x"00",x"0f",x"3f"),
    11 => (x"30",x"18",x"30",x"7f"),
    12 => (x"41",x"00",x"7f",x"7f"),
    13 => (x"1c",x"1c",x"36",x"63"),
    14 => (x"01",x"41",x"63",x"36"),
    15 => (x"7c",x"7c",x"06",x"03"),
    16 => (x"61",x"01",x"03",x"06"),
    17 => (x"47",x"4d",x"59",x"71"),
    18 => (x"00",x"00",x"41",x"43"),
    19 => (x"41",x"7f",x"7f",x"00"),
    20 => (x"01",x"00",x"00",x"41"),
    21 => (x"18",x"0c",x"06",x"03"),
    22 => (x"00",x"40",x"60",x"30"),
    23 => (x"7f",x"41",x"41",x"00"),
    24 => (x"08",x"00",x"00",x"7f"),
    25 => (x"06",x"03",x"06",x"0c"),
    26 => (x"80",x"00",x"08",x"0c"),
    27 => (x"80",x"80",x"80",x"80"),
    28 => (x"00",x"00",x"80",x"80"),
    29 => (x"07",x"03",x"00",x"00"),
    30 => (x"00",x"00",x"00",x"04"),
    31 => (x"54",x"54",x"74",x"20"),
    32 => (x"00",x"00",x"78",x"7c"),
    33 => (x"44",x"44",x"7f",x"7f"),
    34 => (x"00",x"00",x"38",x"7c"),
    35 => (x"44",x"44",x"7c",x"38"),
    36 => (x"00",x"00",x"00",x"44"),
    37 => (x"44",x"44",x"7c",x"38"),
    38 => (x"00",x"00",x"7f",x"7f"),
    39 => (x"54",x"54",x"7c",x"38"),
    40 => (x"00",x"00",x"18",x"5c"),
    41 => (x"05",x"7f",x"7e",x"04"),
    42 => (x"00",x"00",x"00",x"05"),
    43 => (x"a4",x"a4",x"bc",x"18"),
    44 => (x"00",x"00",x"7c",x"fc"),
    45 => (x"04",x"04",x"7f",x"7f"),
    46 => (x"00",x"00",x"78",x"7c"),
    47 => (x"7d",x"3d",x"00",x"00"),
    48 => (x"00",x"00",x"00",x"40"),
    49 => (x"fd",x"80",x"80",x"80"),
    50 => (x"00",x"00",x"00",x"7d"),
    51 => (x"38",x"10",x"7f",x"7f"),
    52 => (x"00",x"00",x"44",x"6c"),
    53 => (x"7f",x"3f",x"00",x"00"),
    54 => (x"7c",x"00",x"00",x"40"),
    55 => (x"0c",x"18",x"0c",x"7c"),
    56 => (x"00",x"00",x"78",x"7c"),
    57 => (x"04",x"04",x"7c",x"7c"),
    58 => (x"00",x"00",x"78",x"7c"),
    59 => (x"44",x"44",x"7c",x"38"),
    60 => (x"00",x"00",x"38",x"7c"),
    61 => (x"24",x"24",x"fc",x"fc"),
    62 => (x"00",x"00",x"18",x"3c"),
    63 => (x"24",x"24",x"3c",x"18"),
    64 => (x"00",x"00",x"fc",x"fc"),
    65 => (x"04",x"04",x"7c",x"7c"),
    66 => (x"00",x"00",x"08",x"0c"),
    67 => (x"54",x"54",x"5c",x"48"),
    68 => (x"00",x"00",x"20",x"74"),
    69 => (x"44",x"7f",x"3f",x"04"),
    70 => (x"00",x"00",x"00",x"44"),
    71 => (x"40",x"40",x"7c",x"3c"),
    72 => (x"00",x"00",x"7c",x"7c"),
    73 => (x"60",x"60",x"3c",x"1c"),
    74 => (x"3c",x"00",x"1c",x"3c"),
    75 => (x"60",x"30",x"60",x"7c"),
    76 => (x"44",x"00",x"3c",x"7c"),
    77 => (x"38",x"10",x"38",x"6c"),
    78 => (x"00",x"00",x"44",x"6c"),
    79 => (x"60",x"e0",x"bc",x"1c"),
    80 => (x"00",x"00",x"1c",x"3c"),
    81 => (x"5c",x"74",x"64",x"44"),
    82 => (x"00",x"00",x"44",x"4c"),
    83 => (x"77",x"3e",x"08",x"08"),
    84 => (x"00",x"00",x"41",x"41"),
    85 => (x"7f",x"7f",x"00",x"00"),
    86 => (x"00",x"00",x"00",x"00"),
    87 => (x"3e",x"77",x"41",x"41"),
    88 => (x"02",x"00",x"08",x"08"),
    89 => (x"02",x"03",x"01",x"01"),
    90 => (x"7f",x"00",x"01",x"02"),
    91 => (x"7f",x"7f",x"7f",x"7f"),
    92 => (x"08",x"00",x"7f",x"7f"),
    93 => (x"3e",x"1c",x"1c",x"08"),
    94 => (x"7f",x"7f",x"7f",x"3e"),
    95 => (x"1c",x"3e",x"3e",x"7f"),
    96 => (x"00",x"08",x"08",x"1c"),
    97 => (x"7c",x"7c",x"18",x"10"),
    98 => (x"00",x"00",x"10",x"18"),
    99 => (x"7c",x"7c",x"30",x"10"),
   100 => (x"10",x"00",x"10",x"30"),
   101 => (x"78",x"60",x"60",x"30"),
   102 => (x"42",x"00",x"06",x"1e"),
   103 => (x"3c",x"18",x"3c",x"66"),
   104 => (x"78",x"00",x"42",x"66"),
   105 => (x"c6",x"c2",x"6a",x"38"),
   106 => (x"60",x"00",x"38",x"6c"),
   107 => (x"00",x"60",x"00",x"00"),
   108 => (x"0e",x"00",x"60",x"00"),
   109 => (x"5d",x"5c",x"5b",x"5e"),
   110 => (x"4c",x"71",x"1e",x"0e"),
   111 => (x"bf",x"fd",x"f0",x"c2"),
   112 => (x"c0",x"4b",x"c0",x"4d"),
   113 => (x"02",x"ab",x"74",x"1e"),
   114 => (x"a6",x"c4",x"87",x"c7"),
   115 => (x"c5",x"78",x"c0",x"48"),
   116 => (x"48",x"a6",x"c4",x"87"),
   117 => (x"66",x"c4",x"78",x"c1"),
   118 => (x"ee",x"49",x"73",x"1e"),
   119 => (x"86",x"c8",x"87",x"df"),
   120 => (x"ef",x"49",x"e0",x"c0"),
   121 => (x"a5",x"c4",x"87",x"ef"),
   122 => (x"f0",x"49",x"6a",x"4a"),
   123 => (x"c6",x"f1",x"87",x"f0"),
   124 => (x"c1",x"85",x"cb",x"87"),
   125 => (x"ab",x"b7",x"c8",x"83"),
   126 => (x"87",x"c7",x"ff",x"04"),
   127 => (x"26",x"4d",x"26",x"26"),
   128 => (x"26",x"4b",x"26",x"4c"),
   129 => (x"4a",x"71",x"1e",x"4f"),
   130 => (x"5a",x"c1",x"f1",x"c2"),
   131 => (x"48",x"c1",x"f1",x"c2"),
   132 => (x"fe",x"49",x"78",x"c7"),
   133 => (x"4f",x"26",x"87",x"dd"),
   134 => (x"71",x"1e",x"73",x"1e"),
   135 => (x"aa",x"b7",x"c0",x"4a"),
   136 => (x"c2",x"87",x"d3",x"03"),
   137 => (x"05",x"bf",x"f2",x"d5"),
   138 => (x"4b",x"c1",x"87",x"c4"),
   139 => (x"4b",x"c0",x"87",x"c2"),
   140 => (x"5b",x"f6",x"d5",x"c2"),
   141 => (x"d5",x"c2",x"87",x"c4"),
   142 => (x"d5",x"c2",x"5a",x"f6"),
   143 => (x"c1",x"4a",x"bf",x"f2"),
   144 => (x"a2",x"c0",x"c1",x"9a"),
   145 => (x"87",x"e8",x"ec",x"49"),
   146 => (x"d5",x"c2",x"48",x"fc"),
   147 => (x"fe",x"78",x"bf",x"f2"),
   148 => (x"71",x"1e",x"87",x"ef"),
   149 => (x"1e",x"66",x"c4",x"4a"),
   150 => (x"e2",x"e6",x"49",x"72"),
   151 => (x"4f",x"26",x"26",x"87"),
   152 => (x"f2",x"d5",x"c2",x"1e"),
   153 => (x"c4",x"e3",x"49",x"bf"),
   154 => (x"f5",x"f0",x"c2",x"87"),
   155 => (x"78",x"bf",x"e8",x"48"),
   156 => (x"48",x"f1",x"f0",x"c2"),
   157 => (x"c2",x"78",x"bf",x"ec"),
   158 => (x"4a",x"bf",x"f5",x"f0"),
   159 => (x"99",x"ff",x"c3",x"49"),
   160 => (x"72",x"2a",x"b7",x"c8"),
   161 => (x"c2",x"b0",x"71",x"48"),
   162 => (x"26",x"58",x"fd",x"f0"),
   163 => (x"5b",x"5e",x"0e",x"4f"),
   164 => (x"71",x"0e",x"5d",x"5c"),
   165 => (x"87",x"c8",x"ff",x"4b"),
   166 => (x"48",x"f0",x"f0",x"c2"),
   167 => (x"49",x"73",x"50",x"c0"),
   168 => (x"70",x"87",x"ea",x"e2"),
   169 => (x"9c",x"c2",x"4c",x"49"),
   170 => (x"cb",x"49",x"ee",x"cb"),
   171 => (x"49",x"70",x"87",x"cc"),
   172 => (x"f0",x"f0",x"c2",x"4d"),
   173 => (x"c1",x"05",x"bf",x"97"),
   174 => (x"66",x"d0",x"87",x"e2"),
   175 => (x"f9",x"f0",x"c2",x"49"),
   176 => (x"d6",x"05",x"99",x"bf"),
   177 => (x"49",x"66",x"d4",x"87"),
   178 => (x"bf",x"f1",x"f0",x"c2"),
   179 => (x"87",x"cb",x"05",x"99"),
   180 => (x"f8",x"e1",x"49",x"73"),
   181 => (x"02",x"98",x"70",x"87"),
   182 => (x"c1",x"87",x"c1",x"c1"),
   183 => (x"87",x"c0",x"fe",x"4c"),
   184 => (x"e1",x"ca",x"49",x"75"),
   185 => (x"02",x"98",x"70",x"87"),
   186 => (x"f0",x"c2",x"87",x"c6"),
   187 => (x"50",x"c1",x"48",x"f0"),
   188 => (x"97",x"f0",x"f0",x"c2"),
   189 => (x"e3",x"c0",x"05",x"bf"),
   190 => (x"f9",x"f0",x"c2",x"87"),
   191 => (x"66",x"d0",x"49",x"bf"),
   192 => (x"d6",x"ff",x"05",x"99"),
   193 => (x"f1",x"f0",x"c2",x"87"),
   194 => (x"66",x"d4",x"49",x"bf"),
   195 => (x"ca",x"ff",x"05",x"99"),
   196 => (x"e0",x"49",x"73",x"87"),
   197 => (x"98",x"70",x"87",x"f7"),
   198 => (x"87",x"ff",x"fe",x"05"),
   199 => (x"dc",x"fb",x"48",x"74"),
   200 => (x"5b",x"5e",x"0e",x"87"),
   201 => (x"f4",x"0e",x"5d",x"5c"),
   202 => (x"4c",x"4d",x"c0",x"86"),
   203 => (x"c4",x"7e",x"bf",x"ec"),
   204 => (x"f0",x"c2",x"48",x"a6"),
   205 => (x"c1",x"78",x"bf",x"fd"),
   206 => (x"c7",x"1e",x"c0",x"1e"),
   207 => (x"87",x"cd",x"fd",x"49"),
   208 => (x"98",x"70",x"86",x"c8"),
   209 => (x"ff",x"87",x"ce",x"02"),
   210 => (x"87",x"cc",x"fb",x"49"),
   211 => (x"ff",x"49",x"da",x"c1"),
   212 => (x"c1",x"87",x"fa",x"df"),
   213 => (x"f0",x"f0",x"c2",x"4d"),
   214 => (x"c3",x"02",x"bf",x"97"),
   215 => (x"87",x"c4",x"d0",x"87"),
   216 => (x"bf",x"f5",x"f0",x"c2"),
   217 => (x"f2",x"d5",x"c2",x"4b"),
   218 => (x"eb",x"c0",x"05",x"bf"),
   219 => (x"49",x"fd",x"c3",x"87"),
   220 => (x"87",x"d9",x"df",x"ff"),
   221 => (x"ff",x"49",x"fa",x"c3"),
   222 => (x"73",x"87",x"d2",x"df"),
   223 => (x"99",x"ff",x"c3",x"49"),
   224 => (x"49",x"c0",x"1e",x"71"),
   225 => (x"73",x"87",x"cb",x"fb"),
   226 => (x"29",x"b7",x"c8",x"49"),
   227 => (x"49",x"c1",x"1e",x"71"),
   228 => (x"c8",x"87",x"ff",x"fa"),
   229 => (x"87",x"c0",x"c6",x"86"),
   230 => (x"bf",x"f9",x"f0",x"c2"),
   231 => (x"dd",x"02",x"9b",x"4b"),
   232 => (x"ee",x"d5",x"c2",x"87"),
   233 => (x"dd",x"c7",x"49",x"bf"),
   234 => (x"05",x"98",x"70",x"87"),
   235 => (x"4b",x"c0",x"87",x"c4"),
   236 => (x"e0",x"c2",x"87",x"d2"),
   237 => (x"87",x"c2",x"c7",x"49"),
   238 => (x"58",x"f2",x"d5",x"c2"),
   239 => (x"d5",x"c2",x"87",x"c6"),
   240 => (x"78",x"c0",x"48",x"ee"),
   241 => (x"99",x"c2",x"49",x"73"),
   242 => (x"c3",x"87",x"ce",x"05"),
   243 => (x"dd",x"ff",x"49",x"eb"),
   244 => (x"49",x"70",x"87",x"fb"),
   245 => (x"c2",x"02",x"99",x"c2"),
   246 => (x"73",x"4c",x"fb",x"87"),
   247 => (x"05",x"99",x"c1",x"49"),
   248 => (x"f4",x"c3",x"87",x"ce"),
   249 => (x"e4",x"dd",x"ff",x"49"),
   250 => (x"c2",x"49",x"70",x"87"),
   251 => (x"87",x"c2",x"02",x"99"),
   252 => (x"49",x"73",x"4c",x"fa"),
   253 => (x"ce",x"05",x"99",x"c8"),
   254 => (x"49",x"f5",x"c3",x"87"),
   255 => (x"87",x"cd",x"dd",x"ff"),
   256 => (x"99",x"c2",x"49",x"70"),
   257 => (x"c2",x"87",x"d5",x"02"),
   258 => (x"02",x"bf",x"c1",x"f1"),
   259 => (x"c1",x"48",x"87",x"ca"),
   260 => (x"c5",x"f1",x"c2",x"88"),
   261 => (x"87",x"c2",x"c0",x"58"),
   262 => (x"4d",x"c1",x"4c",x"ff"),
   263 => (x"99",x"c4",x"49",x"73"),
   264 => (x"c3",x"87",x"ce",x"05"),
   265 => (x"dc",x"ff",x"49",x"f2"),
   266 => (x"49",x"70",x"87",x"e3"),
   267 => (x"dc",x"02",x"99",x"c2"),
   268 => (x"c1",x"f1",x"c2",x"87"),
   269 => (x"c7",x"48",x"7e",x"bf"),
   270 => (x"c0",x"03",x"a8",x"b7"),
   271 => (x"48",x"6e",x"87",x"cb"),
   272 => (x"f1",x"c2",x"80",x"c1"),
   273 => (x"c2",x"c0",x"58",x"c5"),
   274 => (x"c1",x"4c",x"fe",x"87"),
   275 => (x"49",x"fd",x"c3",x"4d"),
   276 => (x"87",x"f9",x"db",x"ff"),
   277 => (x"99",x"c2",x"49",x"70"),
   278 => (x"c2",x"87",x"d5",x"02"),
   279 => (x"02",x"bf",x"c1",x"f1"),
   280 => (x"c2",x"87",x"c9",x"c0"),
   281 => (x"c0",x"48",x"c1",x"f1"),
   282 => (x"87",x"c2",x"c0",x"78"),
   283 => (x"4d",x"c1",x"4c",x"fd"),
   284 => (x"ff",x"49",x"fa",x"c3"),
   285 => (x"70",x"87",x"d6",x"db"),
   286 => (x"02",x"99",x"c2",x"49"),
   287 => (x"c2",x"87",x"d9",x"c0"),
   288 => (x"48",x"bf",x"c1",x"f1"),
   289 => (x"03",x"a8",x"b7",x"c7"),
   290 => (x"c2",x"87",x"c9",x"c0"),
   291 => (x"c7",x"48",x"c1",x"f1"),
   292 => (x"87",x"c2",x"c0",x"78"),
   293 => (x"4d",x"c1",x"4c",x"fc"),
   294 => (x"03",x"ac",x"b7",x"c0"),
   295 => (x"c4",x"87",x"d1",x"c0"),
   296 => (x"d8",x"c1",x"4a",x"66"),
   297 => (x"c0",x"02",x"6a",x"82"),
   298 => (x"4b",x"6a",x"87",x"c6"),
   299 => (x"0f",x"73",x"49",x"74"),
   300 => (x"f0",x"c3",x"1e",x"c0"),
   301 => (x"49",x"da",x"c1",x"1e"),
   302 => (x"c8",x"87",x"d2",x"f7"),
   303 => (x"02",x"98",x"70",x"86"),
   304 => (x"c8",x"87",x"e2",x"c0"),
   305 => (x"f1",x"c2",x"48",x"a6"),
   306 => (x"c8",x"78",x"bf",x"c1"),
   307 => (x"91",x"cb",x"49",x"66"),
   308 => (x"71",x"48",x"66",x"c4"),
   309 => (x"6e",x"7e",x"70",x"80"),
   310 => (x"c8",x"c0",x"02",x"bf"),
   311 => (x"4b",x"bf",x"6e",x"87"),
   312 => (x"73",x"49",x"66",x"c8"),
   313 => (x"02",x"9d",x"75",x"0f"),
   314 => (x"c2",x"87",x"c8",x"c0"),
   315 => (x"49",x"bf",x"c1",x"f1"),
   316 => (x"c2",x"87",x"c0",x"f3"),
   317 => (x"02",x"bf",x"f6",x"d5"),
   318 => (x"49",x"87",x"dd",x"c0"),
   319 => (x"70",x"87",x"c7",x"c2"),
   320 => (x"d3",x"c0",x"02",x"98"),
   321 => (x"c1",x"f1",x"c2",x"87"),
   322 => (x"e6",x"f2",x"49",x"bf"),
   323 => (x"f4",x"49",x"c0",x"87"),
   324 => (x"d5",x"c2",x"87",x"c6"),
   325 => (x"78",x"c0",x"48",x"f6"),
   326 => (x"e0",x"f3",x"8e",x"f4"),
   327 => (x"5b",x"5e",x"0e",x"87"),
   328 => (x"1e",x"0e",x"5d",x"5c"),
   329 => (x"f0",x"c2",x"4c",x"71"),
   330 => (x"c1",x"49",x"bf",x"fd"),
   331 => (x"c1",x"4d",x"a1",x"cd"),
   332 => (x"7e",x"69",x"81",x"d1"),
   333 => (x"cf",x"02",x"9c",x"74"),
   334 => (x"4b",x"a5",x"c4",x"87"),
   335 => (x"f0",x"c2",x"7b",x"74"),
   336 => (x"f2",x"49",x"bf",x"fd"),
   337 => (x"7b",x"6e",x"87",x"ff"),
   338 => (x"c4",x"05",x"9c",x"74"),
   339 => (x"c2",x"4b",x"c0",x"87"),
   340 => (x"73",x"4b",x"c1",x"87"),
   341 => (x"87",x"c0",x"f3",x"49"),
   342 => (x"c7",x"02",x"66",x"d4"),
   343 => (x"87",x"da",x"49",x"87"),
   344 => (x"87",x"c2",x"4a",x"70"),
   345 => (x"d5",x"c2",x"4a",x"c0"),
   346 => (x"f2",x"26",x"5a",x"fa"),
   347 => (x"00",x"00",x"87",x"cf"),
   348 => (x"00",x"00",x"00",x"00"),
   349 => (x"00",x"00",x"00",x"00"),
   350 => (x"71",x"1e",x"00",x"00"),
   351 => (x"bf",x"c8",x"ff",x"4a"),
   352 => (x"48",x"a1",x"72",x"49"),
   353 => (x"ff",x"1e",x"4f",x"26"),
   354 => (x"fe",x"89",x"bf",x"c8"),
   355 => (x"c0",x"c0",x"c0",x"c0"),
   356 => (x"c4",x"01",x"a9",x"c0"),
   357 => (x"c2",x"4a",x"c0",x"87"),
   358 => (x"72",x"4a",x"c1",x"87"),
   359 => (x"0e",x"4f",x"26",x"48"),
   360 => (x"5d",x"5c",x"5b",x"5e"),
   361 => (x"ff",x"4b",x"71",x"0e"),
   362 => (x"66",x"d0",x"4c",x"d4"),
   363 => (x"d6",x"78",x"c0",x"48"),
   364 => (x"d0",x"d8",x"ff",x"49"),
   365 => (x"7c",x"ff",x"c3",x"87"),
   366 => (x"ff",x"c3",x"49",x"6c"),
   367 => (x"49",x"4d",x"71",x"99"),
   368 => (x"c1",x"99",x"f0",x"c3"),
   369 => (x"cb",x"05",x"a9",x"e0"),
   370 => (x"7c",x"ff",x"c3",x"87"),
   371 => (x"98",x"c3",x"48",x"6c"),
   372 => (x"78",x"08",x"66",x"d0"),
   373 => (x"6c",x"7c",x"ff",x"c3"),
   374 => (x"31",x"c8",x"49",x"4a"),
   375 => (x"6c",x"7c",x"ff",x"c3"),
   376 => (x"72",x"b2",x"71",x"4a"),
   377 => (x"c3",x"31",x"c8",x"49"),
   378 => (x"4a",x"6c",x"7c",x"ff"),
   379 => (x"49",x"72",x"b2",x"71"),
   380 => (x"ff",x"c3",x"31",x"c8"),
   381 => (x"71",x"4a",x"6c",x"7c"),
   382 => (x"48",x"d0",x"ff",x"b2"),
   383 => (x"73",x"78",x"e0",x"c0"),
   384 => (x"87",x"c2",x"02",x"9b"),
   385 => (x"48",x"75",x"7b",x"72"),
   386 => (x"4c",x"26",x"4d",x"26"),
   387 => (x"4f",x"26",x"4b",x"26"),
   388 => (x"0e",x"4f",x"26",x"1e"),
   389 => (x"0e",x"5c",x"5b",x"5e"),
   390 => (x"1e",x"76",x"86",x"f8"),
   391 => (x"fd",x"49",x"a6",x"c8"),
   392 => (x"86",x"c4",x"87",x"fd"),
   393 => (x"48",x"6e",x"4b",x"70"),
   394 => (x"c2",x"03",x"a8",x"c2"),
   395 => (x"4a",x"73",x"87",x"f0"),
   396 => (x"c1",x"9a",x"f0",x"c3"),
   397 => (x"c7",x"02",x"aa",x"d0"),
   398 => (x"aa",x"e0",x"c1",x"87"),
   399 => (x"87",x"de",x"c2",x"05"),
   400 => (x"99",x"c8",x"49",x"73"),
   401 => (x"ff",x"87",x"c3",x"02"),
   402 => (x"4c",x"73",x"87",x"c6"),
   403 => (x"ac",x"c2",x"9c",x"c3"),
   404 => (x"87",x"c2",x"c1",x"05"),
   405 => (x"c9",x"49",x"66",x"c4"),
   406 => (x"c4",x"1e",x"71",x"31"),
   407 => (x"92",x"d4",x"4a",x"66"),
   408 => (x"49",x"c5",x"f1",x"c2"),
   409 => (x"cd",x"fe",x"81",x"72"),
   410 => (x"49",x"d8",x"87",x"f6"),
   411 => (x"87",x"d5",x"d5",x"ff"),
   412 => (x"c2",x"1e",x"c0",x"c8"),
   413 => (x"fd",x"49",x"de",x"df"),
   414 => (x"ff",x"87",x"f1",x"e9"),
   415 => (x"e0",x"c0",x"48",x"d0"),
   416 => (x"de",x"df",x"c2",x"78"),
   417 => (x"4a",x"66",x"cc",x"1e"),
   418 => (x"f1",x"c2",x"92",x"d4"),
   419 => (x"81",x"72",x"49",x"c5"),
   420 => (x"87",x"fd",x"cb",x"fe"),
   421 => (x"ac",x"c1",x"86",x"cc"),
   422 => (x"87",x"c2",x"c1",x"05"),
   423 => (x"c9",x"49",x"66",x"c4"),
   424 => (x"c4",x"1e",x"71",x"31"),
   425 => (x"92",x"d4",x"4a",x"66"),
   426 => (x"49",x"c5",x"f1",x"c2"),
   427 => (x"cc",x"fe",x"81",x"72"),
   428 => (x"df",x"c2",x"87",x"ee"),
   429 => (x"66",x"c8",x"1e",x"de"),
   430 => (x"c2",x"92",x"d4",x"4a"),
   431 => (x"72",x"49",x"c5",x"f1"),
   432 => (x"fd",x"c9",x"fe",x"81"),
   433 => (x"ff",x"49",x"d7",x"87"),
   434 => (x"c8",x"87",x"fa",x"d3"),
   435 => (x"df",x"c2",x"1e",x"c0"),
   436 => (x"e7",x"fd",x"49",x"de"),
   437 => (x"86",x"cc",x"87",x"ef"),
   438 => (x"c0",x"48",x"d0",x"ff"),
   439 => (x"8e",x"f8",x"78",x"e0"),
   440 => (x"0e",x"87",x"e7",x"fc"),
   441 => (x"5d",x"5c",x"5b",x"5e"),
   442 => (x"4d",x"71",x"1e",x"0e"),
   443 => (x"d4",x"4c",x"d4",x"ff"),
   444 => (x"c3",x"48",x"7e",x"66"),
   445 => (x"c5",x"06",x"a8",x"b7"),
   446 => (x"c1",x"48",x"c0",x"87"),
   447 => (x"49",x"75",x"87",x"e2"),
   448 => (x"87",x"c2",x"db",x"fe"),
   449 => (x"66",x"c4",x"1e",x"75"),
   450 => (x"c2",x"93",x"d4",x"4b"),
   451 => (x"73",x"83",x"c5",x"f1"),
   452 => (x"d8",x"c5",x"fe",x"49"),
   453 => (x"6b",x"83",x"c8",x"87"),
   454 => (x"48",x"d0",x"ff",x"4b"),
   455 => (x"dd",x"78",x"e1",x"c8"),
   456 => (x"c3",x"49",x"73",x"7c"),
   457 => (x"7c",x"71",x"99",x"ff"),
   458 => (x"b7",x"c8",x"49",x"73"),
   459 => (x"99",x"ff",x"c3",x"29"),
   460 => (x"49",x"73",x"7c",x"71"),
   461 => (x"c3",x"29",x"b7",x"d0"),
   462 => (x"7c",x"71",x"99",x"ff"),
   463 => (x"b7",x"d8",x"49",x"73"),
   464 => (x"c0",x"7c",x"71",x"29"),
   465 => (x"7c",x"7c",x"7c",x"7c"),
   466 => (x"7c",x"7c",x"7c",x"7c"),
   467 => (x"7c",x"7c",x"7c",x"7c"),
   468 => (x"c4",x"78",x"e0",x"c0"),
   469 => (x"49",x"dc",x"1e",x"66"),
   470 => (x"87",x"ce",x"d2",x"ff"),
   471 => (x"48",x"73",x"86",x"c8"),
   472 => (x"87",x"e4",x"fa",x"26"),
   473 => (x"f2",x"de",x"c2",x"1e"),
   474 => (x"b9",x"c1",x"49",x"bf"),
   475 => (x"59",x"f6",x"de",x"c2"),
   476 => (x"c3",x"48",x"d4",x"ff"),
   477 => (x"d0",x"ff",x"78",x"ff"),
   478 => (x"78",x"e1",x"c0",x"48"),
   479 => (x"c1",x"48",x"d4",x"ff"),
   480 => (x"71",x"31",x"c4",x"78"),
   481 => (x"48",x"d0",x"ff",x"78"),
   482 => (x"26",x"78",x"e0",x"c0"),
   483 => (x"de",x"c2",x"1e",x"4f"),
   484 => (x"ec",x"c2",x"1e",x"e6"),
   485 => (x"c3",x"fe",x"49",x"d4"),
   486 => (x"86",x"c4",x"87",x"d3"),
   487 => (x"c3",x"02",x"98",x"70"),
   488 => (x"87",x"c0",x"ff",x"87"),
   489 => (x"35",x"31",x"4f",x"26"),
   490 => (x"20",x"5a",x"48",x"4b"),
   491 => (x"46",x"43",x"20",x"20"),
   492 => (x"00",x"00",x"00",x"47"),
   493 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

