library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f4f1c287",
    12 => x"86c0c64e",
    13 => x"49f4f1c2",
    14 => x"48fcdec2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087dde1",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"4a711e4f",
    50 => x"484966c4",
    51 => x"a6c888c1",
    52 => x"02997158",
    53 => x"481287d4",
    54 => x"7808d4ff",
    55 => x"484966c4",
    56 => x"a6c888c1",
    57 => x"05997158",
    58 => x"4f2687ec",
    59 => x"c44a711e",
    60 => x"c1484966",
    61 => x"58a6c888",
    62 => x"d6029971",
    63 => x"48d4ff87",
    64 => x"6878ffc3",
    65 => x"4966c452",
    66 => x"c888c148",
    67 => x"997158a6",
    68 => x"2687ea05",
    69 => x"1e731e4f",
    70 => x"c34bd4ff",
    71 => x"4a6b7bff",
    72 => x"6b7bffc3",
    73 => x"7232c849",
    74 => x"7bffc3b1",
    75 => x"31c84a6b",
    76 => x"ffc3b271",
    77 => x"c8496b7b",
    78 => x"71b17232",
    79 => x"2687c448",
    80 => x"264c264d",
    81 => x"0e4f264b",
    82 => x"5d5c5b5e",
    83 => x"ff4a710e",
    84 => x"49724cd4",
    85 => x"7199ffc3",
    86 => x"fcdec27c",
    87 => x"87c805bf",
    88 => x"c94866d0",
    89 => x"58a6d430",
    90 => x"d84966d0",
    91 => x"99ffc329",
    92 => x"66d07c71",
    93 => x"c329d049",
    94 => x"7c7199ff",
    95 => x"c84966d0",
    96 => x"99ffc329",
    97 => x"66d07c71",
    98 => x"99ffc349",
    99 => x"49727c71",
   100 => x"ffc329d0",
   101 => x"6c7c7199",
   102 => x"fff0c94b",
   103 => x"abffc34d",
   104 => x"c387d005",
   105 => x"4b6c7cff",
   106 => x"c6028dc1",
   107 => x"abffc387",
   108 => x"7387f002",
   109 => x"87c7fe48",
   110 => x"ff49c01e",
   111 => x"ffc348d4",
   112 => x"c381c178",
   113 => x"04a9b7c8",
   114 => x"4f2687f1",
   115 => x"e71e731e",
   116 => x"dff8c487",
   117 => x"c01ec04b",
   118 => x"f7c1f0ff",
   119 => x"87e7fd49",
   120 => x"a8c186c4",
   121 => x"87eac005",
   122 => x"c348d4ff",
   123 => x"c0c178ff",
   124 => x"c0c0c0c0",
   125 => x"f0e1c01e",
   126 => x"fd49e9c1",
   127 => x"86c487c9",
   128 => x"ca059870",
   129 => x"48d4ff87",
   130 => x"c178ffc3",
   131 => x"fe87cb48",
   132 => x"8bc187e6",
   133 => x"87fdfe05",
   134 => x"e6fc48c0",
   135 => x"1e731e87",
   136 => x"c348d4ff",
   137 => x"4bd378ff",
   138 => x"ffc01ec0",
   139 => x"49c1c1f0",
   140 => x"c487d4fc",
   141 => x"05987086",
   142 => x"d4ff87ca",
   143 => x"78ffc348",
   144 => x"87cb48c1",
   145 => x"c187f1fd",
   146 => x"dbff058b",
   147 => x"fb48c087",
   148 => x"5e0e87f1",
   149 => x"ff0e5c5b",
   150 => x"dbfd4cd4",
   151 => x"1eeac687",
   152 => x"c1f0e1c0",
   153 => x"defb49c8",
   154 => x"c186c487",
   155 => x"87c802a8",
   156 => x"c087eafe",
   157 => x"87e2c148",
   158 => x"7087dafa",
   159 => x"ffffcf49",
   160 => x"a9eac699",
   161 => x"fe87c802",
   162 => x"48c087d3",
   163 => x"c387cbc1",
   164 => x"f1c07cff",
   165 => x"87f4fc4b",
   166 => x"c0029870",
   167 => x"1ec087eb",
   168 => x"c1f0ffc0",
   169 => x"defa49fa",
   170 => x"7086c487",
   171 => x"87d90598",
   172 => x"6c7cffc3",
   173 => x"7cffc349",
   174 => x"c17c7c7c",
   175 => x"c40299c0",
   176 => x"d548c187",
   177 => x"d148c087",
   178 => x"05abc287",
   179 => x"48c087c4",
   180 => x"8bc187c8",
   181 => x"87fdfe05",
   182 => x"e4f948c0",
   183 => x"1e731e87",
   184 => x"48fcdec2",
   185 => x"4bc778c1",
   186 => x"c248d0ff",
   187 => x"87c8fb78",
   188 => x"c348d0ff",
   189 => x"c01ec078",
   190 => x"c0c1d0e5",
   191 => x"87c7f949",
   192 => x"a8c186c4",
   193 => x"4b87c105",
   194 => x"c505abc2",
   195 => x"c048c087",
   196 => x"8bc187f9",
   197 => x"87d0ff05",
   198 => x"c287f7fc",
   199 => x"7058c0df",
   200 => x"87cd0598",
   201 => x"ffc01ec1",
   202 => x"49d0c1f0",
   203 => x"c487d8f8",
   204 => x"48d4ff86",
   205 => x"c478ffc3",
   206 => x"dfc287de",
   207 => x"d0ff58c4",
   208 => x"ff78c248",
   209 => x"ffc348d4",
   210 => x"f748c178",
   211 => x"5e0e87f5",
   212 => x"0e5d5c5b",
   213 => x"ffc34a71",
   214 => x"4cd4ff4d",
   215 => x"d0ff7c75",
   216 => x"78c3c448",
   217 => x"1e727c75",
   218 => x"c1f0ffc0",
   219 => x"d6f749d8",
   220 => x"7086c487",
   221 => x"87c50298",
   222 => x"f0c048c1",
   223 => x"c37c7587",
   224 => x"c0c87cfe",
   225 => x"4966d41e",
   226 => x"c487faf4",
   227 => x"757c7586",
   228 => x"d87c757c",
   229 => x"754be0da",
   230 => x"99496c7c",
   231 => x"c187c505",
   232 => x"87f3058b",
   233 => x"d0ff7c75",
   234 => x"c078c248",
   235 => x"87cff648",
   236 => x"5c5b5e0e",
   237 => x"4b710e5d",
   238 => x"eec54cc0",
   239 => x"ff4adfcd",
   240 => x"ffc348d4",
   241 => x"c3496878",
   242 => x"c005a9fe",
   243 => x"4d7087fd",
   244 => x"cc029b73",
   245 => x"1e66d087",
   246 => x"cff44973",
   247 => x"d686c487",
   248 => x"48d0ff87",
   249 => x"c378d1c4",
   250 => x"66d07dff",
   251 => x"d488c148",
   252 => x"987058a6",
   253 => x"ff87f005",
   254 => x"ffc348d4",
   255 => x"9b737878",
   256 => x"ff87c505",
   257 => x"78d048d0",
   258 => x"c14c4ac1",
   259 => x"eefe058a",
   260 => x"f4487487",
   261 => x"731e87e9",
   262 => x"c04a711e",
   263 => x"48d4ff4b",
   264 => x"ff78ffc3",
   265 => x"c3c448d0",
   266 => x"48d4ff78",
   267 => x"7278ffc3",
   268 => x"f0ffc01e",
   269 => x"f449d1c1",
   270 => x"86c487cd",
   271 => x"d2059870",
   272 => x"1ec0c887",
   273 => x"fd4966cc",
   274 => x"86c487e6",
   275 => x"d0ff4b70",
   276 => x"7378c248",
   277 => x"87ebf348",
   278 => x"5c5b5e0e",
   279 => x"1ec00e5d",
   280 => x"c1f0ffc0",
   281 => x"def349c9",
   282 => x"c21ed287",
   283 => x"fc49c4df",
   284 => x"86c887fe",
   285 => x"84c14cc0",
   286 => x"04acb7d2",
   287 => x"dfc287f8",
   288 => x"49bf97c4",
   289 => x"c199c0c3",
   290 => x"c005a9c0",
   291 => x"dfc287e7",
   292 => x"49bf97cb",
   293 => x"dfc231d0",
   294 => x"4abf97cc",
   295 => x"b17232c8",
   296 => x"97cddfc2",
   297 => x"71b14abf",
   298 => x"ffffcf4c",
   299 => x"84c19cff",
   300 => x"e7c134ca",
   301 => x"cddfc287",
   302 => x"c149bf97",
   303 => x"c299c631",
   304 => x"bf97cedf",
   305 => x"2ab7c74a",
   306 => x"dfc2b172",
   307 => x"4abf97c9",
   308 => x"c29dcf4d",
   309 => x"bf97cadf",
   310 => x"ca9ac34a",
   311 => x"cbdfc232",
   312 => x"c24bbf97",
   313 => x"c2b27333",
   314 => x"bf97ccdf",
   315 => x"9bc0c34b",
   316 => x"732bb7c6",
   317 => x"c181c2b2",
   318 => x"70307148",
   319 => x"7548c149",
   320 => x"724d7030",
   321 => x"7184c14c",
   322 => x"b7c0c894",
   323 => x"87cc06ad",
   324 => x"2db734c1",
   325 => x"adb7c0c8",
   326 => x"87f4ff01",
   327 => x"def04874",
   328 => x"5b5e0e87",
   329 => x"f80e5d5c",
   330 => x"eae7c286",
   331 => x"c278c048",
   332 => x"c01ee2df",
   333 => x"87defb49",
   334 => x"987086c4",
   335 => x"c087c505",
   336 => x"87cec948",
   337 => x"7ec14dc0",
   338 => x"bfc0f3c0",
   339 => x"d8e0c249",
   340 => x"4bc8714a",
   341 => x"7087d3ec",
   342 => x"87c20598",
   343 => x"f2c07ec0",
   344 => x"c249bffc",
   345 => x"714af4e0",
   346 => x"fdeb4bc8",
   347 => x"05987087",
   348 => x"7ec087c2",
   349 => x"fdc0026e",
   350 => x"e8e6c287",
   351 => x"e7c24dbf",
   352 => x"7ebf9fe0",
   353 => x"ead6c548",
   354 => x"87c705a8",
   355 => x"bfe8e6c2",
   356 => x"6e87ce4d",
   357 => x"d5e9ca48",
   358 => x"87c502a8",
   359 => x"f1c748c0",
   360 => x"e2dfc287",
   361 => x"f949751e",
   362 => x"86c487ec",
   363 => x"c5059870",
   364 => x"c748c087",
   365 => x"f2c087dc",
   366 => x"c249bffc",
   367 => x"714af4e0",
   368 => x"e5ea4bc8",
   369 => x"05987087",
   370 => x"e7c287c8",
   371 => x"78c148ea",
   372 => x"f3c087da",
   373 => x"c249bfc0",
   374 => x"714ad8e0",
   375 => x"c9ea4bc8",
   376 => x"02987087",
   377 => x"c087c5c0",
   378 => x"87e6c648",
   379 => x"97e0e7c2",
   380 => x"d5c149bf",
   381 => x"cdc005a9",
   382 => x"e1e7c287",
   383 => x"c249bf97",
   384 => x"c002a9ea",
   385 => x"48c087c5",
   386 => x"c287c7c6",
   387 => x"bf97e2df",
   388 => x"e9c3487e",
   389 => x"cec002a8",
   390 => x"c3486e87",
   391 => x"c002a8eb",
   392 => x"48c087c5",
   393 => x"c287ebc5",
   394 => x"bf97eddf",
   395 => x"c0059949",
   396 => x"dfc287cc",
   397 => x"49bf97ee",
   398 => x"c002a9c2",
   399 => x"48c087c5",
   400 => x"c287cfc5",
   401 => x"bf97efdf",
   402 => x"e6e7c248",
   403 => x"484c7058",
   404 => x"e7c288c1",
   405 => x"dfc258ea",
   406 => x"49bf97f0",
   407 => x"dfc28175",
   408 => x"4abf97f1",
   409 => x"a17232c8",
   410 => x"f7ebc27e",
   411 => x"c2786e48",
   412 => x"bf97f2df",
   413 => x"58a6c848",
   414 => x"bfeae7c2",
   415 => x"87d4c202",
   416 => x"bffcf2c0",
   417 => x"f4e0c249",
   418 => x"4bc8714a",
   419 => x"7087dbe7",
   420 => x"c5c00298",
   421 => x"c348c087",
   422 => x"e7c287f8",
   423 => x"c24cbfe2",
   424 => x"c25ccbec",
   425 => x"bf97c7e0",
   426 => x"c231c849",
   427 => x"bf97c6e0",
   428 => x"c249a14a",
   429 => x"bf97c8e0",
   430 => x"7232d04a",
   431 => x"e0c249a1",
   432 => x"4abf97c9",
   433 => x"a17232d8",
   434 => x"9166c449",
   435 => x"bff7ebc2",
   436 => x"ffebc281",
   437 => x"cfe0c259",
   438 => x"c84abf97",
   439 => x"cee0c232",
   440 => x"a24bbf97",
   441 => x"d0e0c24a",
   442 => x"d04bbf97",
   443 => x"4aa27333",
   444 => x"97d1e0c2",
   445 => x"9bcf4bbf",
   446 => x"a27333d8",
   447 => x"c3ecc24a",
   448 => x"ffebc25a",
   449 => x"8ac24abf",
   450 => x"ecc29274",
   451 => x"a17248c3",
   452 => x"87cac178",
   453 => x"97f4dfc2",
   454 => x"31c849bf",
   455 => x"97f3dfc2",
   456 => x"49a14abf",
   457 => x"59f2e7c2",
   458 => x"bfeee7c2",
   459 => x"c731c549",
   460 => x"29c981ff",
   461 => x"59cbecc2",
   462 => x"97f9dfc2",
   463 => x"32c84abf",
   464 => x"97f8dfc2",
   465 => x"4aa24bbf",
   466 => x"6e9266c4",
   467 => x"c7ecc282",
   468 => x"ffebc25a",
   469 => x"c278c048",
   470 => x"7248fbeb",
   471 => x"ecc278a1",
   472 => x"ebc248cb",
   473 => x"c278bfff",
   474 => x"c248cfec",
   475 => x"78bfc3ec",
   476 => x"bfeae7c2",
   477 => x"87c9c002",
   478 => x"30c44874",
   479 => x"c9c07e70",
   480 => x"c7ecc287",
   481 => x"30c448bf",
   482 => x"e7c27e70",
   483 => x"786e48ee",
   484 => x"8ef848c1",
   485 => x"4c264d26",
   486 => x"4f264b26",
   487 => x"5c5b5e0e",
   488 => x"4a710e5d",
   489 => x"bfeae7c2",
   490 => x"7287cb02",
   491 => x"722bc74b",
   492 => x"9cffc14c",
   493 => x"4b7287c9",
   494 => x"4c722bc8",
   495 => x"c29cffc3",
   496 => x"83bff7eb",
   497 => x"bff8f2c0",
   498 => x"87d902ab",
   499 => x"5bfcf2c0",
   500 => x"1ee2dfc2",
   501 => x"fdf04973",
   502 => x"7086c487",
   503 => x"87c50598",
   504 => x"e6c048c0",
   505 => x"eae7c287",
   506 => x"87d202bf",
   507 => x"91c44974",
   508 => x"81e2dfc2",
   509 => x"ffcf4d69",
   510 => x"9dffffff",
   511 => x"497487cb",
   512 => x"dfc291c2",
   513 => x"699f81e2",
   514 => x"fe48754d",
   515 => x"5e0e87c6",
   516 => x"0e5d5c5b",
   517 => x"c04d711e",
   518 => x"ca49c11e",
   519 => x"86c487ff",
   520 => x"029c4c70",
   521 => x"c287c0c1",
   522 => x"754af2e7",
   523 => x"87dfe049",
   524 => x"c0029870",
   525 => x"4a7487f1",
   526 => x"4bcb4975",
   527 => x"7087c5e1",
   528 => x"e2c00298",
   529 => x"741ec087",
   530 => x"87c7029c",
   531 => x"c048a6c4",
   532 => x"c487c578",
   533 => x"78c148a6",
   534 => x"c94966c4",
   535 => x"86c487ff",
   536 => x"059c4c70",
   537 => x"7487c0ff",
   538 => x"e7fc2648",
   539 => x"5b5e0e87",
   540 => x"1e0e5d5c",
   541 => x"059b4b71",
   542 => x"48c087c5",
   543 => x"c887e5c1",
   544 => x"7dc04da3",
   545 => x"c70266d4",
   546 => x"9766d487",
   547 => x"87c505bf",
   548 => x"cfc148c0",
   549 => x"4966d487",
   550 => x"7087f3fd",
   551 => x"c1029c4c",
   552 => x"a4dc87c0",
   553 => x"da7d6949",
   554 => x"a3c449a4",
   555 => x"7a699f4a",
   556 => x"bfeae7c2",
   557 => x"d487d202",
   558 => x"699f49a4",
   559 => x"ffffc049",
   560 => x"d0487199",
   561 => x"c27e7030",
   562 => x"6e7ec087",
   563 => x"806a4849",
   564 => x"7bc07a70",
   565 => x"6a49a3cc",
   566 => x"49a3d079",
   567 => x"48c179c0",
   568 => x"48c087c2",
   569 => x"87ecfa26",
   570 => x"5c5b5e0e",
   571 => x"4c710e5d",
   572 => x"cac1029c",
   573 => x"49a4c887",
   574 => x"c2c10269",
   575 => x"4a66d087",
   576 => x"d482496c",
   577 => x"66d05aa6",
   578 => x"e7c2b94d",
   579 => x"ff4abfe6",
   580 => x"719972ba",
   581 => x"e4c00299",
   582 => x"4ba4c487",
   583 => x"fbf9496b",
   584 => x"c27b7087",
   585 => x"49bfe2e7",
   586 => x"7c71816c",
   587 => x"e7c2b975",
   588 => x"ff4abfe6",
   589 => x"719972ba",
   590 => x"dcff0599",
   591 => x"f97c7587",
   592 => x"731e87d2",
   593 => x"9b4b711e",
   594 => x"c887c702",
   595 => x"056949a3",
   596 => x"48c087c5",
   597 => x"c287f7c0",
   598 => x"4abffbeb",
   599 => x"6949a3c4",
   600 => x"c289c249",
   601 => x"91bfe2e7",
   602 => x"c24aa271",
   603 => x"49bfe6e7",
   604 => x"a271996b",
   605 => x"fcf2c04a",
   606 => x"1e66c85a",
   607 => x"d5ea4972",
   608 => x"7086c487",
   609 => x"87c40598",
   610 => x"87c248c0",
   611 => x"c7f848c1",
   612 => x"1e731e87",
   613 => x"029b4b71",
   614 => x"a3c887c7",
   615 => x"c5056949",
   616 => x"c048c087",
   617 => x"ebc287f7",
   618 => x"c44abffb",
   619 => x"496949a3",
   620 => x"e7c289c2",
   621 => x"7191bfe2",
   622 => x"e7c24aa2",
   623 => x"6b49bfe6",
   624 => x"4aa27199",
   625 => x"5afcf2c0",
   626 => x"721e66c8",
   627 => x"87fee549",
   628 => x"987086c4",
   629 => x"c087c405",
   630 => x"c187c248",
   631 => x"87f8f648",
   632 => x"5c5b5e0e",
   633 => x"711e0e5d",
   634 => x"4c66d44b",
   635 => x"9b732cc9",
   636 => x"87cfc102",
   637 => x"6949a3c8",
   638 => x"87c7c102",
   639 => x"d44da3d0",
   640 => x"e7c27d66",
   641 => x"ff49bfe6",
   642 => x"994a6bb9",
   643 => x"03ac717e",
   644 => x"7bc087cd",
   645 => x"4aa3cc7d",
   646 => x"6a49a3c4",
   647 => x"7287c279",
   648 => x"029c748c",
   649 => x"1e4987dd",
   650 => x"fbfa4973",
   651 => x"d486c487",
   652 => x"ffc74966",
   653 => x"87cb0299",
   654 => x"1ee2dfc2",
   655 => x"c1fc4973",
   656 => x"2686c487",
   657 => x"1e87cdf5",
   658 => x"4b711e73",
   659 => x"e4c0029b",
   660 => x"cfecc287",
   661 => x"c24a735b",
   662 => x"e2e7c28a",
   663 => x"c29249bf",
   664 => x"48bffbeb",
   665 => x"ecc28072",
   666 => x"487158d3",
   667 => x"e7c230c4",
   668 => x"edc058f2",
   669 => x"cbecc287",
   670 => x"ffebc248",
   671 => x"ecc278bf",
   672 => x"ecc248cf",
   673 => x"c278bfc3",
   674 => x"02bfeae7",
   675 => x"e7c287c9",
   676 => x"c449bfe2",
   677 => x"c287c731",
   678 => x"49bfc7ec",
   679 => x"e7c231c4",
   680 => x"f3f359f2",
   681 => x"5b5e0e87",
   682 => x"4a710e5c",
   683 => x"9a724bc0",
   684 => x"87e1c002",
   685 => x"9f49a2da",
   686 => x"e7c24b69",
   687 => x"cf02bfea",
   688 => x"49a2d487",
   689 => x"4c49699f",
   690 => x"9cffffc0",
   691 => x"87c234d0",
   692 => x"49744cc0",
   693 => x"fd4973b3",
   694 => x"f9f287ed",
   695 => x"5b5e0e87",
   696 => x"f40e5d5c",
   697 => x"c04a7186",
   698 => x"029a727e",
   699 => x"dfc287d8",
   700 => x"78c048de",
   701 => x"48d6dfc2",
   702 => x"bfcfecc2",
   703 => x"dadfc278",
   704 => x"cbecc248",
   705 => x"e7c278bf",
   706 => x"50c048ff",
   707 => x"bfeee7c2",
   708 => x"dedfc249",
   709 => x"aa714abf",
   710 => x"87c9c403",
   711 => x"99cf4972",
   712 => x"87e9c005",
   713 => x"48f8f2c0",
   714 => x"bfd6dfc2",
   715 => x"e2dfc278",
   716 => x"d6dfc21e",
   717 => x"dfc249bf",
   718 => x"a1c148d6",
   719 => x"d5e37178",
   720 => x"c086c487",
   721 => x"c248f4f2",
   722 => x"cc78e2df",
   723 => x"f4f2c087",
   724 => x"e0c048bf",
   725 => x"f8f2c080",
   726 => x"dedfc258",
   727 => x"80c148bf",
   728 => x"58e2dfc2",
   729 => x"000cb427",
   730 => x"bf97bf00",
   731 => x"c2029d4d",
   732 => x"e5c387e3",
   733 => x"dcc202ad",
   734 => x"f4f2c087",
   735 => x"a3cb4bbf",
   736 => x"cf4c1149",
   737 => x"d2c105ac",
   738 => x"df497587",
   739 => x"cd89c199",
   740 => x"f2e7c291",
   741 => x"4aa3c181",
   742 => x"a3c35112",
   743 => x"c551124a",
   744 => x"51124aa3",
   745 => x"124aa3c7",
   746 => x"4aa3c951",
   747 => x"a3ce5112",
   748 => x"d051124a",
   749 => x"51124aa3",
   750 => x"124aa3d2",
   751 => x"4aa3d451",
   752 => x"a3d65112",
   753 => x"d851124a",
   754 => x"51124aa3",
   755 => x"124aa3dc",
   756 => x"4aa3de51",
   757 => x"7ec15112",
   758 => x"7487fac0",
   759 => x"0599c849",
   760 => x"7487ebc0",
   761 => x"0599d049",
   762 => x"66dc87d1",
   763 => x"87cbc002",
   764 => x"66dc4973",
   765 => x"0298700f",
   766 => x"6e87d3c0",
   767 => x"87c6c005",
   768 => x"48f2e7c2",
   769 => x"f2c050c0",
   770 => x"c248bff4",
   771 => x"e7c287e1",
   772 => x"50c048ff",
   773 => x"eee7c27e",
   774 => x"dfc249bf",
   775 => x"714abfde",
   776 => x"f7fb04aa",
   777 => x"cfecc287",
   778 => x"c8c005bf",
   779 => x"eae7c287",
   780 => x"f8c102bf",
   781 => x"dadfc287",
   782 => x"dfed49bf",
   783 => x"c2497087",
   784 => x"c459dedf",
   785 => x"dfc248a6",
   786 => x"c278bfda",
   787 => x"02bfeae7",
   788 => x"c487d8c0",
   789 => x"ffcf4966",
   790 => x"99f8ffff",
   791 => x"c5c002a9",
   792 => x"c04cc087",
   793 => x"4cc187e1",
   794 => x"c487dcc0",
   795 => x"ffcf4966",
   796 => x"02a999f8",
   797 => x"c887c8c0",
   798 => x"78c048a6",
   799 => x"c887c5c0",
   800 => x"78c148a6",
   801 => x"744c66c8",
   802 => x"e0c0059c",
   803 => x"4966c487",
   804 => x"e7c289c2",
   805 => x"914abfe2",
   806 => x"bffbebc2",
   807 => x"d6dfc24a",
   808 => x"78a17248",
   809 => x"48dedfc2",
   810 => x"dff978c0",
   811 => x"f448c087",
   812 => x"87e0eb8e",
   813 => x"00000000",
   814 => x"ffffffff",
   815 => x"00000cc4",
   816 => x"00000ccd",
   817 => x"33544146",
   818 => x"20202032",
   819 => x"54414600",
   820 => x"20203631",
   821 => x"ff1e0020",
   822 => x"ffc348d4",
   823 => x"26486878",
   824 => x"d4ff1e4f",
   825 => x"78ffc348",
   826 => x"c848d0ff",
   827 => x"d4ff78e1",
   828 => x"c278d448",
   829 => x"ff48d3ec",
   830 => x"2650bfd4",
   831 => x"d0ff1e4f",
   832 => x"78e0c048",
   833 => x"ff1e4f26",
   834 => x"497087cc",
   835 => x"87c60299",
   836 => x"05a9fbc0",
   837 => x"487187f1",
   838 => x"5e0e4f26",
   839 => x"710e5c5b",
   840 => x"fe4cc04b",
   841 => x"497087f0",
   842 => x"f9c00299",
   843 => x"a9ecc087",
   844 => x"87f2c002",
   845 => x"02a9fbc0",
   846 => x"cc87ebc0",
   847 => x"03acb766",
   848 => x"66d087c7",
   849 => x"7187c202",
   850 => x"02997153",
   851 => x"84c187c2",
   852 => x"7087c3fe",
   853 => x"cd029949",
   854 => x"a9ecc087",
   855 => x"c087c702",
   856 => x"ff05a9fb",
   857 => x"66d087d5",
   858 => x"c087c302",
   859 => x"ecc07b97",
   860 => x"87c405a9",
   861 => x"87c54a74",
   862 => x"0ac04a74",
   863 => x"c248728a",
   864 => x"264d2687",
   865 => x"264b264c",
   866 => x"c9fd1e4f",
   867 => x"c0497087",
   868 => x"04a9b7f0",
   869 => x"f9c087ca",
   870 => x"c301a9b7",
   871 => x"89f0c087",
   872 => x"a9b7c1c1",
   873 => x"c187ca04",
   874 => x"01a9b7da",
   875 => x"f7c087c3",
   876 => x"b7e1c189",
   877 => x"87ca04a9",
   878 => x"a9b7fac1",
   879 => x"c087c301",
   880 => x"487189fd",
   881 => x"5e0e4f26",
   882 => x"710e5c5b",
   883 => x"4cd4ff4a",
   884 => x"eac04972",
   885 => x"9b4b7087",
   886 => x"c187c202",
   887 => x"48d0ff8b",
   888 => x"c178c5c8",
   889 => x"49737cd5",
   890 => x"e2c131c6",
   891 => x"4abf97fe",
   892 => x"70b07148",
   893 => x"48d0ff7c",
   894 => x"487378c4",
   895 => x"0e87c4fe",
   896 => x"5d5c5b5e",
   897 => x"7186f80e",
   898 => x"fb7ec04c",
   899 => x"4bc087d3",
   900 => x"97ecfac0",
   901 => x"a9c049bf",
   902 => x"fb87cf04",
   903 => x"83c187e8",
   904 => x"97ecfac0",
   905 => x"06ab49bf",
   906 => x"fac087f1",
   907 => x"02bf97ec",
   908 => x"e1fa87cf",
   909 => x"99497087",
   910 => x"c087c602",
   911 => x"f105a9ec",
   912 => x"fa4bc087",
   913 => x"4d7087d0",
   914 => x"c887cbfa",
   915 => x"c5fa58a6",
   916 => x"c14a7087",
   917 => x"49a4c883",
   918 => x"ad496997",
   919 => x"c087c702",
   920 => x"c005adff",
   921 => x"a4c987e7",
   922 => x"49699749",
   923 => x"02a966c4",
   924 => x"c04887c7",
   925 => x"d405a8ff",
   926 => x"49a4ca87",
   927 => x"aa496997",
   928 => x"c087c602",
   929 => x"c405aaff",
   930 => x"d07ec187",
   931 => x"adecc087",
   932 => x"c087c602",
   933 => x"c405adfb",
   934 => x"c14bc087",
   935 => x"fe026e7e",
   936 => x"d8f987e1",
   937 => x"f8487387",
   938 => x"87d5fb8e",
   939 => x"5b5e0e00",
   940 => x"1e0e5d5c",
   941 => x"d4ff4d71",
   942 => x"c21e754b",
   943 => x"e649d8ec",
   944 => x"86c487eb",
   945 => x"c3029870",
   946 => x"ecc287d8",
   947 => x"754cbfe0",
   948 => x"87f2fb49",
   949 => x"c848d0ff",
   950 => x"d6c178c5",
   951 => x"754ac07b",
   952 => x"7b1149a2",
   953 => x"b7cb82c1",
   954 => x"87f304aa",
   955 => x"ffc34acc",
   956 => x"c082c17b",
   957 => x"04aab7e0",
   958 => x"d0ff87f4",
   959 => x"c378c448",
   960 => x"c5c87bff",
   961 => x"7bd3c178",
   962 => x"78c47bc1",
   963 => x"c1029c74",
   964 => x"dfc287ff",
   965 => x"c0c87ee2",
   966 => x"b7c08c4d",
   967 => x"87c603ac",
   968 => x"4da4c0c8",
   969 => x"c0c84cc0",
   970 => x"87dc05ad",
   971 => x"97d3ecc2",
   972 => x"99d049bf",
   973 => x"c087d102",
   974 => x"d8ecc21e",
   975 => x"87c2e849",
   976 => x"497086c4",
   977 => x"87eec04a",
   978 => x"1ee2dfc2",
   979 => x"49d8ecc2",
   980 => x"c487efe7",
   981 => x"4a497086",
   982 => x"c848d0ff",
   983 => x"d4c178c5",
   984 => x"bf976e7b",
   985 => x"c1486e7b",
   986 => x"c17e7080",
   987 => x"f0ff058d",
   988 => x"48d0ff87",
   989 => x"9a7278c4",
   990 => x"c087c505",
   991 => x"87e4c048",
   992 => x"ecc21ec1",
   993 => x"dfe549d8",
   994 => x"7486c487",
   995 => x"c1fe059c",
   996 => x"48d0ff87",
   997 => x"c178c5c8",
   998 => x"7bc07bd3",
   999 => x"48c178c4",
  1000 => x"48c087c2",
  1001 => x"264d2626",
  1002 => x"264b264c",
  1003 => x"5b5e0e4f",
  1004 => x"1e0e5d5c",
  1005 => x"4cc04b71",
  1006 => x"c004ab4d",
  1007 => x"f7c087e8",
  1008 => x"9d751eff",
  1009 => x"c087c402",
  1010 => x"c187c24a",
  1011 => x"ec49724a",
  1012 => x"86c487cb",
  1013 => x"84c17e70",
  1014 => x"87c2056e",
  1015 => x"85c14c73",
  1016 => x"ff06ac73",
  1017 => x"486e87d8",
  1018 => x"87f9fe26",
  1019 => x"5c5b5e0e",
  1020 => x"cc4b710e",
  1021 => x"87d80266",
  1022 => x"8cf0c04c",
  1023 => x"7487d802",
  1024 => x"028ac14a",
  1025 => x"028a87d1",
  1026 => x"028a87cd",
  1027 => x"87d987c9",
  1028 => x"d8fa4973",
  1029 => x"7487d287",
  1030 => x"c149c01e",
  1031 => x"7487c8db",
  1032 => x"c149731e",
  1033 => x"c887c0db",
  1034 => x"87fbfd86",
  1035 => x"5c5b5e0e",
  1036 => x"711e0e5d",
  1037 => x"91de494c",
  1038 => x"4dc0edc2",
  1039 => x"6d978571",
  1040 => x"87dcc102",
  1041 => x"bfececc2",
  1042 => x"7282744a",
  1043 => x"87ddfd49",
  1044 => x"026e7e70",
  1045 => x"c287f2c0",
  1046 => x"6e4bf4ec",
  1047 => x"ff49cb4a",
  1048 => x"7487c5c1",
  1049 => x"c193cb4b",
  1050 => x"c483cee3",
  1051 => x"e4c2c183",
  1052 => x"c149747b",
  1053 => x"7587c0c5",
  1054 => x"ffe2c17b",
  1055 => x"1e49bf97",
  1056 => x"49f4ecc2",
  1057 => x"c487e5fd",
  1058 => x"c1497486",
  1059 => x"c087e8c4",
  1060 => x"c7c6c149",
  1061 => x"d4ecc287",
  1062 => x"c178c048",
  1063 => x"87ffdc49",
  1064 => x"87c1fc26",
  1065 => x"64616f4c",
  1066 => x"2e676e69",
  1067 => x"0e002e2e",
  1068 => x"0e5c5b5e",
  1069 => x"c24a4b71",
  1070 => x"82bfecec",
  1071 => x"ecfb4972",
  1072 => x"9c4c7087",
  1073 => x"4987c402",
  1074 => x"c287dae7",
  1075 => x"c048ecec",
  1076 => x"dc49c178",
  1077 => x"cefb87c9",
  1078 => x"5b5e0e87",
  1079 => x"f40e5d5c",
  1080 => x"e2dfc286",
  1081 => x"c44cc04d",
  1082 => x"78c048a6",
  1083 => x"bfececc2",
  1084 => x"06a9c049",
  1085 => x"c287c1c1",
  1086 => x"9848e2df",
  1087 => x"87f8c002",
  1088 => x"1efff7c0",
  1089 => x"c70266c8",
  1090 => x"48a6c487",
  1091 => x"87c578c0",
  1092 => x"c148a6c4",
  1093 => x"4966c478",
  1094 => x"c487c2e7",
  1095 => x"c14d7086",
  1096 => x"4866c484",
  1097 => x"a6c880c1",
  1098 => x"ececc258",
  1099 => x"03ac49bf",
  1100 => x"9d7587c6",
  1101 => x"87c8ff05",
  1102 => x"9d754cc0",
  1103 => x"87e0c302",
  1104 => x"1efff7c0",
  1105 => x"c70266c8",
  1106 => x"48a6cc87",
  1107 => x"87c578c0",
  1108 => x"c148a6cc",
  1109 => x"4966cc78",
  1110 => x"c487c2e6",
  1111 => x"6e7e7086",
  1112 => x"87e9c202",
  1113 => x"81cb496e",
  1114 => x"d0496997",
  1115 => x"d6c10299",
  1116 => x"efc2c187",
  1117 => x"cb49744a",
  1118 => x"cee3c191",
  1119 => x"c8797281",
  1120 => x"51ffc381",
  1121 => x"91de4974",
  1122 => x"4dc0edc2",
  1123 => x"c1c28571",
  1124 => x"a5c17d97",
  1125 => x"51e0c049",
  1126 => x"97f2e7c2",
  1127 => x"87d202bf",
  1128 => x"a5c284c1",
  1129 => x"f2e7c24b",
  1130 => x"fe49db4a",
  1131 => x"c187f9fb",
  1132 => x"a5cd87db",
  1133 => x"c151c049",
  1134 => x"4ba5c284",
  1135 => x"49cb4a6e",
  1136 => x"87e4fbfe",
  1137 => x"c187c6c1",
  1138 => x"744aecc0",
  1139 => x"c191cb49",
  1140 => x"7281cee3",
  1141 => x"f2e7c279",
  1142 => x"d802bf97",
  1143 => x"de497487",
  1144 => x"c284c191",
  1145 => x"714bc0ed",
  1146 => x"f2e7c283",
  1147 => x"fe49dd4a",
  1148 => x"d887f5fa",
  1149 => x"de4b7487",
  1150 => x"c0edc293",
  1151 => x"49a3cb83",
  1152 => x"84c151c0",
  1153 => x"cb4a6e73",
  1154 => x"dbfafe49",
  1155 => x"4866c487",
  1156 => x"a6c880c1",
  1157 => x"03acc758",
  1158 => x"6e87c5c0",
  1159 => x"87e0fc05",
  1160 => x"8ef44874",
  1161 => x"1e87fef5",
  1162 => x"4b711e73",
  1163 => x"c191cb49",
  1164 => x"c881cee3",
  1165 => x"e2c14aa1",
  1166 => x"501248fe",
  1167 => x"c04aa1c9",
  1168 => x"1248ecfa",
  1169 => x"c181ca50",
  1170 => x"1148ffe2",
  1171 => x"ffe2c150",
  1172 => x"1e49bf97",
  1173 => x"d3f649c0",
  1174 => x"d4ecc287",
  1175 => x"c178de48",
  1176 => x"87fbd549",
  1177 => x"87c1f526",
  1178 => x"494a711e",
  1179 => x"e3c191cb",
  1180 => x"81c881ce",
  1181 => x"ecc24811",
  1182 => x"ecc258d8",
  1183 => x"78c048ec",
  1184 => x"dad549c1",
  1185 => x"1e4f2687",
  1186 => x"fec049c0",
  1187 => x"4f2687ce",
  1188 => x"0299711e",
  1189 => x"e4c187d2",
  1190 => x"50c048e3",
  1191 => x"c9c180f7",
  1192 => x"e3c140e8",
  1193 => x"87ce78c7",
  1194 => x"48dfe4c1",
  1195 => x"78c0e3c1",
  1196 => x"cac180fc",
  1197 => x"4f2678c7",
  1198 => x"5c5b5e0e",
  1199 => x"4a4c710e",
  1200 => x"e3c192cb",
  1201 => x"a2c882ce",
  1202 => x"4ba2c949",
  1203 => x"1e4b6b97",
  1204 => x"1e496997",
  1205 => x"491282ca",
  1206 => x"87c7e7c0",
  1207 => x"fed349c0",
  1208 => x"c0497487",
  1209 => x"f887d0fb",
  1210 => x"87fbf28e",
  1211 => x"711e731e",
  1212 => x"c3ff494b",
  1213 => x"fe497387",
  1214 => x"ecf287fe",
  1215 => x"1e731e87",
  1216 => x"a3c64b71",
  1217 => x"87db024a",
  1218 => x"d6028ac1",
  1219 => x"c1028a87",
  1220 => x"028a87da",
  1221 => x"8a87fcc0",
  1222 => x"87e1c002",
  1223 => x"87cb028a",
  1224 => x"c787dbc1",
  1225 => x"87c0fd49",
  1226 => x"c287dec1",
  1227 => x"02bfecec",
  1228 => x"4887cbc1",
  1229 => x"ecc288c1",
  1230 => x"c1c158f0",
  1231 => x"f0ecc287",
  1232 => x"f9c002bf",
  1233 => x"ececc287",
  1234 => x"80c148bf",
  1235 => x"58f0ecc2",
  1236 => x"c287ebc0",
  1237 => x"49bfecec",
  1238 => x"ecc289c6",
  1239 => x"b7c059f0",
  1240 => x"87da03a9",
  1241 => x"48ececc2",
  1242 => x"87d278c0",
  1243 => x"bff0ecc2",
  1244 => x"c287cb02",
  1245 => x"48bfecec",
  1246 => x"ecc280c6",
  1247 => x"49c058f0",
  1248 => x"7387dcd1",
  1249 => x"eef8c049",
  1250 => x"87ddf087",
  1251 => x"5c5b5e0e",
  1252 => x"cc4c710e",
  1253 => x"4b741e66",
  1254 => x"e3c193cb",
  1255 => x"a3c483ce",
  1256 => x"fe496a4a",
  1257 => x"c187d1f4",
  1258 => x"c87be7c8",
  1259 => x"66d449a3",
  1260 => x"49a3c951",
  1261 => x"ca5166d8",
  1262 => x"66dc49a3",
  1263 => x"e6ef2651",
  1264 => x"5b5e0e87",
  1265 => x"ff0e5d5c",
  1266 => x"a6d886d0",
  1267 => x"48a6c459",
  1268 => x"80c478c0",
  1269 => x"7866c4c1",
  1270 => x"78c180c4",
  1271 => x"78c180c4",
  1272 => x"48f0ecc2",
  1273 => x"ecc278c1",
  1274 => x"de48bfd4",
  1275 => x"87cb05a8",
  1276 => x"7087e6f3",
  1277 => x"59a6c849",
  1278 => x"e387ecce",
  1279 => x"c5e487e3",
  1280 => x"87d2e387",
  1281 => x"fbc04c70",
  1282 => x"d0c102ac",
  1283 => x"0566d487",
  1284 => x"c087c2c1",
  1285 => x"1ec11e1e",
  1286 => x"1ec1e5c1",
  1287 => x"ebfd49c0",
  1288 => x"66d0c187",
  1289 => x"6a82c44a",
  1290 => x"7481c749",
  1291 => x"d81ec151",
  1292 => x"c8496a1e",
  1293 => x"87e2e381",
  1294 => x"c4c186d8",
  1295 => x"a8c04866",
  1296 => x"c487c701",
  1297 => x"78c148a6",
  1298 => x"c4c187ce",
  1299 => x"88c14866",
  1300 => x"c358a6cc",
  1301 => x"87eee287",
  1302 => x"c248a6cc",
  1303 => x"029c7478",
  1304 => x"c487c0cd",
  1305 => x"c8c14866",
  1306 => x"cc03a866",
  1307 => x"a6d887f5",
  1308 => x"c478c048",
  1309 => x"e178c080",
  1310 => x"4c7087dc",
  1311 => x"05acd0c1",
  1312 => x"dc87d8c2",
  1313 => x"c0e47e66",
  1314 => x"c0497087",
  1315 => x"e159a6e0",
  1316 => x"4c7087c4",
  1317 => x"05acecc0",
  1318 => x"c487ebc1",
  1319 => x"91cb4966",
  1320 => x"8166c0c1",
  1321 => x"6a4aa1c4",
  1322 => x"4aa1c84d",
  1323 => x"c15266dc",
  1324 => x"e079e8c9",
  1325 => x"4c7087e0",
  1326 => x"87d8029c",
  1327 => x"02acfbc0",
  1328 => x"557487d2",
  1329 => x"7087cfe0",
  1330 => x"c7029c4c",
  1331 => x"acfbc087",
  1332 => x"87eeff05",
  1333 => x"c255e0c0",
  1334 => x"97c055c1",
  1335 => x"4966d47d",
  1336 => x"db05a96e",
  1337 => x"4866c487",
  1338 => x"04a866c8",
  1339 => x"66c487ca",
  1340 => x"c880c148",
  1341 => x"87c858a6",
  1342 => x"c14866c8",
  1343 => x"58a6cc88",
  1344 => x"87d2dfff",
  1345 => x"d0c14c70",
  1346 => x"87c805ac",
  1347 => x"c14866d0",
  1348 => x"58a6d480",
  1349 => x"02acd0c1",
  1350 => x"c087e8fd",
  1351 => x"d448a6e0",
  1352 => x"66dc7866",
  1353 => x"66e0c048",
  1354 => x"c8c905a8",
  1355 => x"a6e4c087",
  1356 => x"7e78c048",
  1357 => x"fbc04874",
  1358 => x"a6ecc088",
  1359 => x"02987058",
  1360 => x"4887cdc8",
  1361 => x"ecc088cb",
  1362 => x"987058a6",
  1363 => x"87d2c102",
  1364 => x"c088c948",
  1365 => x"7058a6ec",
  1366 => x"dbc30298",
  1367 => x"88c44887",
  1368 => x"58a6ecc0",
  1369 => x"d0029870",
  1370 => x"88c14887",
  1371 => x"58a6ecc0",
  1372 => x"c3029870",
  1373 => x"d1c787c2",
  1374 => x"48a6d887",
  1375 => x"ff78f0c0",
  1376 => x"7087d3dd",
  1377 => x"acecc04c",
  1378 => x"87c3c002",
  1379 => x"c05ca6dc",
  1380 => x"cd02acec",
  1381 => x"fddcff87",
  1382 => x"c04c7087",
  1383 => x"ff05acec",
  1384 => x"ecc087f3",
  1385 => x"c4c002ac",
  1386 => x"e9dcff87",
  1387 => x"1e66d887",
  1388 => x"1e4966d4",
  1389 => x"1e4966d4",
  1390 => x"1ec1e5c1",
  1391 => x"f74966d4",
  1392 => x"1ec087ca",
  1393 => x"66dc1eca",
  1394 => x"c191cb49",
  1395 => x"d88166d8",
  1396 => x"a1c448a6",
  1397 => x"bf66d878",
  1398 => x"fddcff49",
  1399 => x"c086d887",
  1400 => x"c106a8b7",
  1401 => x"1ec187c5",
  1402 => x"66c81ede",
  1403 => x"dcff49bf",
  1404 => x"86c887e8",
  1405 => x"c0484970",
  1406 => x"a6dc8808",
  1407 => x"a8b7c058",
  1408 => x"87e7c006",
  1409 => x"dd4866d8",
  1410 => x"de03a8b7",
  1411 => x"49bf6e87",
  1412 => x"c08166d8",
  1413 => x"66d851e0",
  1414 => x"6e81c149",
  1415 => x"c1c281bf",
  1416 => x"4966d851",
  1417 => x"bf6e81c2",
  1418 => x"cc51c081",
  1419 => x"80c14866",
  1420 => x"c158a6d0",
  1421 => x"87d8c47e",
  1422 => x"87cdddff",
  1423 => x"ff58a6dc",
  1424 => x"c087c6dd",
  1425 => x"c058a6ec",
  1426 => x"c005a8ec",
  1427 => x"e8c087ca",
  1428 => x"66d848a6",
  1429 => x"87c4c078",
  1430 => x"87fad9ff",
  1431 => x"cb4966c4",
  1432 => x"66c0c191",
  1433 => x"70807148",
  1434 => x"c8496e7e",
  1435 => x"ca4a6e81",
  1436 => x"5266d882",
  1437 => x"4a66e8c0",
  1438 => x"66d882c1",
  1439 => x"7248c18a",
  1440 => x"c14a7030",
  1441 => x"7997728a",
  1442 => x"1e496997",
  1443 => x"d74966dc",
  1444 => x"86c487d3",
  1445 => x"58a6f0c0",
  1446 => x"81c4496e",
  1447 => x"e0c04d69",
  1448 => x"66dc4866",
  1449 => x"c8c002a8",
  1450 => x"48a6d887",
  1451 => x"c5c078c0",
  1452 => x"48a6d887",
  1453 => x"66d878c1",
  1454 => x"1ee0c01e",
  1455 => x"d9ff4975",
  1456 => x"86c887d8",
  1457 => x"b7c04c70",
  1458 => x"d4c106ac",
  1459 => x"c0857487",
  1460 => x"897449e0",
  1461 => x"dfc14b75",
  1462 => x"fe714adc",
  1463 => x"c287c9e7",
  1464 => x"66e4c085",
  1465 => x"c080c148",
  1466 => x"c058a6e8",
  1467 => x"c14966ec",
  1468 => x"02a97081",
  1469 => x"d887c8c0",
  1470 => x"78c048a6",
  1471 => x"d887c5c0",
  1472 => x"78c148a6",
  1473 => x"c21e66d8",
  1474 => x"e0c049a4",
  1475 => x"70887148",
  1476 => x"49751e49",
  1477 => x"87c2d8ff",
  1478 => x"b7c086c8",
  1479 => x"c0ff01a8",
  1480 => x"66e4c087",
  1481 => x"87d1c002",
  1482 => x"81c9496e",
  1483 => x"5166e4c0",
  1484 => x"cac1486e",
  1485 => x"ccc078f8",
  1486 => x"c9496e87",
  1487 => x"6e51c281",
  1488 => x"eccbc148",
  1489 => x"c07ec178",
  1490 => x"d6ff87c6",
  1491 => x"4c7087f8",
  1492 => x"f5c0026e",
  1493 => x"4866c487",
  1494 => x"04a866c8",
  1495 => x"c487cbc0",
  1496 => x"80c14866",
  1497 => x"c058a6c8",
  1498 => x"66c887e0",
  1499 => x"cc88c148",
  1500 => x"d5c058a6",
  1501 => x"acc6c187",
  1502 => x"87c8c005",
  1503 => x"c14866cc",
  1504 => x"58a6d080",
  1505 => x"87fed5ff",
  1506 => x"66d04c70",
  1507 => x"d480c148",
  1508 => x"9c7458a6",
  1509 => x"87cbc002",
  1510 => x"c14866c4",
  1511 => x"04a866c8",
  1512 => x"ff87cbf3",
  1513 => x"c487d6d5",
  1514 => x"a8c74866",
  1515 => x"87e5c003",
  1516 => x"48f0ecc2",
  1517 => x"66c478c0",
  1518 => x"c191cb49",
  1519 => x"c48166c0",
  1520 => x"4a6a4aa1",
  1521 => x"c47952c0",
  1522 => x"80c14866",
  1523 => x"c758a6c8",
  1524 => x"dbff04a8",
  1525 => x"8ed0ff87",
  1526 => x"87c9dfff",
  1527 => x"1e00203a",
  1528 => x"4b711e73",
  1529 => x"87c6029b",
  1530 => x"48ececc2",
  1531 => x"1ec778c0",
  1532 => x"bfececc2",
  1533 => x"e3c11e49",
  1534 => x"ecc21ece",
  1535 => x"ee49bfd4",
  1536 => x"86cc87ff",
  1537 => x"bfd4ecc2",
  1538 => x"87c4ea49",
  1539 => x"c8029b73",
  1540 => x"cee3c187",
  1541 => x"f0e7c049",
  1542 => x"ccdeff87",
  1543 => x"e2c11e87",
  1544 => x"50c048fe",
  1545 => x"bff1e4c1",
  1546 => x"c0daff49",
  1547 => x"2648c087",
  1548 => x"ebc71e4f",
  1549 => x"fe49c187",
  1550 => x"eafe87e5",
  1551 => x"987087df",
  1552 => x"fe87cd02",
  1553 => x"7087daf3",
  1554 => x"87c40298",
  1555 => x"87c24ac1",
  1556 => x"9a724ac0",
  1557 => x"c087ce05",
  1558 => x"c5e2c11e",
  1559 => x"c0f3c049",
  1560 => x"fe86c487",
  1561 => x"e8fcc087",
  1562 => x"c11ec087",
  1563 => x"c049d0e2",
  1564 => x"c087eef2",
  1565 => x"87e5fe1e",
  1566 => x"f2c04970",
  1567 => x"dec387e3",
  1568 => x"268ef887",
  1569 => x"2044534f",
  1570 => x"6c696166",
  1571 => x"002e6465",
  1572 => x"746f6f42",
  1573 => x"2e676e69",
  1574 => x"1e002e2e",
  1575 => x"87c5eac0",
  1576 => x"87f3f5c0",
  1577 => x"4f2687f6",
  1578 => x"ececc21e",
  1579 => x"c278c048",
  1580 => x"c048d4ec",
  1581 => x"87f9fd78",
  1582 => x"48c087e1",
  1583 => x"00004f26",
  1584 => x"78452080",
  1585 => x"80007469",
  1586 => x"63614220",
  1587 => x"1268006b",
  1588 => x"2b400000",
  1589 => x"00000000",
  1590 => x"00126800",
  1591 => x"002b5e00",
  1592 => x"00000000",
  1593 => x"00001268",
  1594 => x"00002b7c",
  1595 => x"68000000",
  1596 => x"9a000012",
  1597 => x"0000002b",
  1598 => x"12680000",
  1599 => x"2bb80000",
  1600 => x"00000000",
  1601 => x"00126800",
  1602 => x"002bd600",
  1603 => x"00000000",
  1604 => x"00001268",
  1605 => x"00002bf4",
  1606 => x"68000000",
  1607 => x"00000012",
  1608 => x"00000000",
  1609 => x"12fd0000",
  1610 => x"00000000",
  1611 => x"00000000",
  1612 => x"00193500",
  1613 => x"34364300",
  1614 => x"20202020",
  1615 => x"4d4f5220",
  1616 => x"616f4c00",
  1617 => x"2e2a2064",
  1618 => x"f0fe1e00",
  1619 => x"cd78c048",
  1620 => x"26097909",
  1621 => x"fe1e1e4f",
  1622 => x"487ebff0",
  1623 => x"1e4f2626",
  1624 => x"c148f0fe",
  1625 => x"1e4f2678",
  1626 => x"c048f0fe",
  1627 => x"1e4f2678",
  1628 => x"52c04a71",
  1629 => x"0e4f2652",
  1630 => x"5d5c5b5e",
  1631 => x"7186f40e",
  1632 => x"7e6d974d",
  1633 => x"974ca5c1",
  1634 => x"a6c8486c",
  1635 => x"c4486e58",
  1636 => x"c505a866",
  1637 => x"c048ff87",
  1638 => x"caff87e6",
  1639 => x"49a5c287",
  1640 => x"714b6c97",
  1641 => x"6b974ba3",
  1642 => x"7e6c974b",
  1643 => x"80c1486e",
  1644 => x"c758a6c8",
  1645 => x"58a6cc98",
  1646 => x"fe7c9770",
  1647 => x"487387e1",
  1648 => x"4d268ef4",
  1649 => x"4b264c26",
  1650 => x"5e0e4f26",
  1651 => x"f40e5c5b",
  1652 => x"d84c7186",
  1653 => x"ffc34a66",
  1654 => x"4ba4c29a",
  1655 => x"73496c97",
  1656 => x"517249a1",
  1657 => x"6e7e6c97",
  1658 => x"c880c148",
  1659 => x"98c758a6",
  1660 => x"7058a6cc",
  1661 => x"ff8ef454",
  1662 => x"1e1e87ca",
  1663 => x"e087e8fd",
  1664 => x"c0494abf",
  1665 => x"0299c0e0",
  1666 => x"1e7287cb",
  1667 => x"49d2f0c2",
  1668 => x"c487f7fe",
  1669 => x"87fdfc86",
  1670 => x"c2fd7e70",
  1671 => x"4f262687",
  1672 => x"d2f0c21e",
  1673 => x"87c7fd49",
  1674 => x"49fae7c1",
  1675 => x"c487dafc",
  1676 => x"4f2687c8",
  1677 => x"48d0ff1e",
  1678 => x"ff78e1c8",
  1679 => x"78c548d4",
  1680 => x"c30266c4",
  1681 => x"78e0c387",
  1682 => x"c60266c8",
  1683 => x"48d4ff87",
  1684 => x"ff78f0c3",
  1685 => x"787148d4",
  1686 => x"c848d0ff",
  1687 => x"e0c078e1",
  1688 => x"0e4f2678",
  1689 => x"0e5c5b5e",
  1690 => x"f0c24c71",
  1691 => x"c6fc49d2",
  1692 => x"c04a7087",
  1693 => x"c204aab7",
  1694 => x"e0c387e3",
  1695 => x"87c905aa",
  1696 => x"48edecc1",
  1697 => x"d4c278c1",
  1698 => x"aaf0c387",
  1699 => x"c187c905",
  1700 => x"c148e9ec",
  1701 => x"87f5c178",
  1702 => x"bfedecc1",
  1703 => x"7287c702",
  1704 => x"b3c0c24b",
  1705 => x"4b7287c2",
  1706 => x"d1059c74",
  1707 => x"e9ecc187",
  1708 => x"ecc11ebf",
  1709 => x"721ebfed",
  1710 => x"87f8fd49",
  1711 => x"ecc186c8",
  1712 => x"c002bfe9",
  1713 => x"497387e0",
  1714 => x"9129b7c4",
  1715 => x"81c9eec1",
  1716 => x"9acf4a73",
  1717 => x"48c192c2",
  1718 => x"4a703072",
  1719 => x"4872baff",
  1720 => x"79709869",
  1721 => x"497387db",
  1722 => x"9129b7c4",
  1723 => x"81c9eec1",
  1724 => x"9acf4a73",
  1725 => x"48c392c2",
  1726 => x"4a703072",
  1727 => x"70b06948",
  1728 => x"edecc179",
  1729 => x"c178c048",
  1730 => x"c048e9ec",
  1731 => x"d2f0c278",
  1732 => x"87e3f949",
  1733 => x"b7c04a70",
  1734 => x"ddfd03aa",
  1735 => x"c248c087",
  1736 => x"264d2687",
  1737 => x"264b264c",
  1738 => x"0000004f",
  1739 => x"00000000",
  1740 => x"4a711e00",
  1741 => x"87ebfc49",
  1742 => x"c01e4f26",
  1743 => x"c449724a",
  1744 => x"c9eec191",
  1745 => x"c179c081",
  1746 => x"aab7d082",
  1747 => x"2687ee04",
  1748 => x"5b5e0e4f",
  1749 => x"710e5d5c",
  1750 => x"87cbf84d",
  1751 => x"b7c44a75",
  1752 => x"eec1922a",
  1753 => x"4c7582c9",
  1754 => x"94c29ccf",
  1755 => x"744b496a",
  1756 => x"c29bc32b",
  1757 => x"70307448",
  1758 => x"74bcff4c",
  1759 => x"70987148",
  1760 => x"87dbf77a",
  1761 => x"d8fe4873",
  1762 => x"00000087",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"d0ff1e00",
  1779 => x"78e1c848",
  1780 => x"d4ff4871",
  1781 => x"4f267808",
  1782 => x"48d0ff1e",
  1783 => x"7178e1c8",
  1784 => x"08d4ff48",
  1785 => x"4866c478",
  1786 => x"7808d4ff",
  1787 => x"711e4f26",
  1788 => x"4966c44a",
  1789 => x"ff49721e",
  1790 => x"d0ff87de",
  1791 => x"78e0c048",
  1792 => x"1e4f2626",
  1793 => x"4b711e73",
  1794 => x"1e4966c8",
  1795 => x"e0c14a73",
  1796 => x"d9ff49a2",
  1797 => x"87c42687",
  1798 => x"4c264d26",
  1799 => x"4f264b26",
  1800 => x"4ad4ff1e",
  1801 => x"ff7affc3",
  1802 => x"e1c848d0",
  1803 => x"c27ade78",
  1804 => x"7abfdcf0",
  1805 => x"28c84849",
  1806 => x"48717a70",
  1807 => x"7a7028d0",
  1808 => x"28d84871",
  1809 => x"f0c27a70",
  1810 => x"497abfe0",
  1811 => x"7028c848",
  1812 => x"d048717a",
  1813 => x"717a7028",
  1814 => x"7028d848",
  1815 => x"48d0ff7a",
  1816 => x"2678e0c0",
  1817 => x"1e731e4f",
  1818 => x"f0c24a71",
  1819 => x"724bbfdc",
  1820 => x"aae0c02b",
  1821 => x"7287ce04",
  1822 => x"89e0c049",
  1823 => x"bfe0f0c2",
  1824 => x"cf2b714b",
  1825 => x"49e0c087",
  1826 => x"f0c28972",
  1827 => x"7148bfe0",
  1828 => x"b3497030",
  1829 => x"739b66c8",
  1830 => x"2687c448",
  1831 => x"264c264d",
  1832 => x"0e4f264b",
  1833 => x"5d5c5b5e",
  1834 => x"7186ec0e",
  1835 => x"dcf0c24b",
  1836 => x"734c7ebf",
  1837 => x"abe0c02c",
  1838 => x"87e0c004",
  1839 => x"c048a6c4",
  1840 => x"c0497378",
  1841 => x"4a7189e0",
  1842 => x"4866e4c0",
  1843 => x"a6cc3072",
  1844 => x"e0f0c258",
  1845 => x"714c4dbf",
  1846 => x"87e4c02c",
  1847 => x"e4c04973",
  1848 => x"30714866",
  1849 => x"c058a6c8",
  1850 => x"897349e0",
  1851 => x"4866e4c0",
  1852 => x"a6cc2871",
  1853 => x"e0f0c258",
  1854 => x"71484dbf",
  1855 => x"b4497030",
  1856 => x"9c66e4c0",
  1857 => x"e8c084c1",
  1858 => x"c204ac66",
  1859 => x"c04cc087",
  1860 => x"d304abe0",
  1861 => x"48a6cc87",
  1862 => x"497378c0",
  1863 => x"7489e0c0",
  1864 => x"d4307148",
  1865 => x"87d558a6",
  1866 => x"48744973",
  1867 => x"a6d03071",
  1868 => x"49e0c058",
  1869 => x"48748973",
  1870 => x"a6d42871",
  1871 => x"4a66c458",
  1872 => x"9a6ebaff",
  1873 => x"ff4966c8",
  1874 => x"729975b9",
  1875 => x"b066cc48",
  1876 => x"58e0f0c2",
  1877 => x"66d04871",
  1878 => x"e4f0c2b0",
  1879 => x"87c0fb58",
  1880 => x"f6fc8eec",
  1881 => x"d0ff1e87",
  1882 => x"78c9c848",
  1883 => x"d4ff4871",
  1884 => x"4f267808",
  1885 => x"494a711e",
  1886 => x"d0ff87eb",
  1887 => x"2678c848",
  1888 => x"1e731e4f",
  1889 => x"f0c24b71",
  1890 => x"c302bff0",
  1891 => x"87ebc287",
  1892 => x"c848d0ff",
  1893 => x"497378c9",
  1894 => x"ffb1e0c0",
  1895 => x"787148d4",
  1896 => x"48e4f0c2",
  1897 => x"66c878c0",
  1898 => x"c387c502",
  1899 => x"87c249ff",
  1900 => x"f0c249c0",
  1901 => x"66cc59ec",
  1902 => x"c587c602",
  1903 => x"c44ad5d5",
  1904 => x"ffffcf87",
  1905 => x"f0f0c24a",
  1906 => x"f0f0c25a",
  1907 => x"c478c148",
  1908 => x"264d2687",
  1909 => x"264b264c",
  1910 => x"5b5e0e4f",
  1911 => x"710e5d5c",
  1912 => x"ecf0c24a",
  1913 => x"9a724cbf",
  1914 => x"4987cb02",
  1915 => x"f5c191c8",
  1916 => x"83714bf7",
  1917 => x"f9c187c4",
  1918 => x"4dc04bf7",
  1919 => x"99744913",
  1920 => x"bfe8f0c2",
  1921 => x"48d4ffb9",
  1922 => x"b7c17871",
  1923 => x"b7c8852c",
  1924 => x"87e804ad",
  1925 => x"bfe4f0c2",
  1926 => x"c280c848",
  1927 => x"fe58e8f0",
  1928 => x"731e87ef",
  1929 => x"134b711e",
  1930 => x"cb029a4a",
  1931 => x"fe497287",
  1932 => x"4a1387e7",
  1933 => x"87f5059a",
  1934 => x"1e87dafe",
  1935 => x"bfe4f0c2",
  1936 => x"e4f0c249",
  1937 => x"78a1c148",
  1938 => x"a9b7c0c4",
  1939 => x"ff87db03",
  1940 => x"f0c248d4",
  1941 => x"c278bfe8",
  1942 => x"49bfe4f0",
  1943 => x"48e4f0c2",
  1944 => x"c478a1c1",
  1945 => x"04a9b7c0",
  1946 => x"d0ff87e5",
  1947 => x"c278c848",
  1948 => x"c048f0f0",
  1949 => x"004f2678",
  1950 => x"00000000",
  1951 => x"00000000",
  1952 => x"5f5f0000",
  1953 => x"00000000",
  1954 => x"03000303",
  1955 => x"14000003",
  1956 => x"7f147f7f",
  1957 => x"0000147f",
  1958 => x"6b6b2e24",
  1959 => x"4c00123a",
  1960 => x"6c18366a",
  1961 => x"30003256",
  1962 => x"77594f7e",
  1963 => x"0040683a",
  1964 => x"03070400",
  1965 => x"00000000",
  1966 => x"633e1c00",
  1967 => x"00000041",
  1968 => x"3e634100",
  1969 => x"0800001c",
  1970 => x"1c1c3e2a",
  1971 => x"00082a3e",
  1972 => x"3e3e0808",
  1973 => x"00000808",
  1974 => x"60e08000",
  1975 => x"00000000",
  1976 => x"08080808",
  1977 => x"00000808",
  1978 => x"60600000",
  1979 => x"40000000",
  1980 => x"0c183060",
  1981 => x"00010306",
  1982 => x"4d597f3e",
  1983 => x"00003e7f",
  1984 => x"7f7f0604",
  1985 => x"00000000",
  1986 => x"59716342",
  1987 => x"0000464f",
  1988 => x"49496322",
  1989 => x"1800367f",
  1990 => x"7f13161c",
  1991 => x"0000107f",
  1992 => x"45456727",
  1993 => x"0000397d",
  1994 => x"494b7e3c",
  1995 => x"00003079",
  1996 => x"79710101",
  1997 => x"0000070f",
  1998 => x"49497f36",
  1999 => x"0000367f",
  2000 => x"69494f06",
  2001 => x"00001e3f",
  2002 => x"66660000",
  2003 => x"00000000",
  2004 => x"66e68000",
  2005 => x"00000000",
  2006 => x"14140808",
  2007 => x"00002222",
  2008 => x"14141414",
  2009 => x"00001414",
  2010 => x"14142222",
  2011 => x"00000808",
  2012 => x"59510302",
  2013 => x"3e00060f",
  2014 => x"555d417f",
  2015 => x"00001e1f",
  2016 => x"09097f7e",
  2017 => x"00007e7f",
  2018 => x"49497f7f",
  2019 => x"0000367f",
  2020 => x"41633e1c",
  2021 => x"00004141",
  2022 => x"63417f7f",
  2023 => x"00001c3e",
  2024 => x"49497f7f",
  2025 => x"00004141",
  2026 => x"09097f7f",
  2027 => x"00000101",
  2028 => x"49417f3e",
  2029 => x"00007a7b",
  2030 => x"08087f7f",
  2031 => x"00007f7f",
  2032 => x"7f7f4100",
  2033 => x"00000041",
  2034 => x"40406020",
  2035 => x"7f003f7f",
  2036 => x"361c087f",
  2037 => x"00004163",
  2038 => x"40407f7f",
  2039 => x"7f004040",
  2040 => x"060c067f",
  2041 => x"7f007f7f",
  2042 => x"180c067f",
  2043 => x"00007f7f",
  2044 => x"41417f3e",
  2045 => x"00003e7f",
  2046 => x"09097f7f",
  2047 => x"3e00060f",
  2048 => x"7f61417f",
  2049 => x"0000407e",
  2050 => x"19097f7f",
  2051 => x"0000667f",
  2052 => x"594d6f26",
  2053 => x"0000327b",
  2054 => x"7f7f0101",
  2055 => x"00000101",
  2056 => x"40407f3f",
  2057 => x"00003f7f",
  2058 => x"70703f0f",
  2059 => x"7f000f3f",
  2060 => x"3018307f",
  2061 => x"41007f7f",
  2062 => x"1c1c3663",
  2063 => x"01416336",
  2064 => x"7c7c0603",
  2065 => x"61010306",
  2066 => x"474d5971",
  2067 => x"00004143",
  2068 => x"417f7f00",
  2069 => x"01000041",
  2070 => x"180c0603",
  2071 => x"00406030",
  2072 => x"7f414100",
  2073 => x"0800007f",
  2074 => x"0603060c",
  2075 => x"8000080c",
  2076 => x"80808080",
  2077 => x"00008080",
  2078 => x"07030000",
  2079 => x"00000004",
  2080 => x"54547420",
  2081 => x"0000787c",
  2082 => x"44447f7f",
  2083 => x"0000387c",
  2084 => x"44447c38",
  2085 => x"00000044",
  2086 => x"44447c38",
  2087 => x"00007f7f",
  2088 => x"54547c38",
  2089 => x"0000185c",
  2090 => x"057f7e04",
  2091 => x"00000005",
  2092 => x"a4a4bc18",
  2093 => x"00007cfc",
  2094 => x"04047f7f",
  2095 => x"0000787c",
  2096 => x"7d3d0000",
  2097 => x"00000040",
  2098 => x"fd808080",
  2099 => x"0000007d",
  2100 => x"38107f7f",
  2101 => x"0000446c",
  2102 => x"7f3f0000",
  2103 => x"7c000040",
  2104 => x"0c180c7c",
  2105 => x"0000787c",
  2106 => x"04047c7c",
  2107 => x"0000787c",
  2108 => x"44447c38",
  2109 => x"0000387c",
  2110 => x"2424fcfc",
  2111 => x"0000183c",
  2112 => x"24243c18",
  2113 => x"0000fcfc",
  2114 => x"04047c7c",
  2115 => x"0000080c",
  2116 => x"54545c48",
  2117 => x"00002074",
  2118 => x"447f3f04",
  2119 => x"00000044",
  2120 => x"40407c3c",
  2121 => x"00007c7c",
  2122 => x"60603c1c",
  2123 => x"3c001c3c",
  2124 => x"6030607c",
  2125 => x"44003c7c",
  2126 => x"3810386c",
  2127 => x"0000446c",
  2128 => x"60e0bc1c",
  2129 => x"00001c3c",
  2130 => x"5c746444",
  2131 => x"0000444c",
  2132 => x"773e0808",
  2133 => x"00004141",
  2134 => x"7f7f0000",
  2135 => x"00000000",
  2136 => x"3e774141",
  2137 => x"02000808",
  2138 => x"02030101",
  2139 => x"7f000102",
  2140 => x"7f7f7f7f",
  2141 => x"08007f7f",
  2142 => x"3e1c1c08",
  2143 => x"7f7f7f3e",
  2144 => x"1c3e3e7f",
  2145 => x"0008081c",
  2146 => x"7c7c1810",
  2147 => x"00001018",
  2148 => x"7c7c3010",
  2149 => x"10001030",
  2150 => x"78606030",
  2151 => x"4200061e",
  2152 => x"3c183c66",
  2153 => x"78004266",
  2154 => x"c6c26a38",
  2155 => x"6000386c",
  2156 => x"00600000",
  2157 => x"0e006000",
  2158 => x"5d5c5b5e",
  2159 => x"4c711e0e",
  2160 => x"bfc1f1c2",
  2161 => x"c04bc04d",
  2162 => x"02ab741e",
  2163 => x"a6c487c7",
  2164 => x"c578c048",
  2165 => x"48a6c487",
  2166 => x"66c478c1",
  2167 => x"ee49731e",
  2168 => x"86c887df",
  2169 => x"ef49e0c0",
  2170 => x"a5c487ef",
  2171 => x"f0496a4a",
  2172 => x"c6f187f0",
  2173 => x"c185cb87",
  2174 => x"abb7c883",
  2175 => x"87c7ff04",
  2176 => x"264d2626",
  2177 => x"264b264c",
  2178 => x"4a711e4f",
  2179 => x"5ac5f1c2",
  2180 => x"48c5f1c2",
  2181 => x"fe4978c7",
  2182 => x"4f2687dd",
  2183 => x"711e731e",
  2184 => x"aab7c04a",
  2185 => x"c287d303",
  2186 => x"05bff6d5",
  2187 => x"4bc187c4",
  2188 => x"4bc087c2",
  2189 => x"5bfad5c2",
  2190 => x"d5c287c4",
  2191 => x"d5c25afa",
  2192 => x"c14abff6",
  2193 => x"a2c0c19a",
  2194 => x"87e8ec49",
  2195 => x"d5c248fc",
  2196 => x"fe78bff6",
  2197 => x"711e87ef",
  2198 => x"1e66c44a",
  2199 => x"e2e64972",
  2200 => x"4f262687",
  2201 => x"f6d5c21e",
  2202 => x"c4e349bf",
  2203 => x"f9f0c287",
  2204 => x"78bfe848",
  2205 => x"48f5f0c2",
  2206 => x"c278bfec",
  2207 => x"4abff9f0",
  2208 => x"99ffc349",
  2209 => x"722ab7c8",
  2210 => x"c2b07148",
  2211 => x"2658c1f1",
  2212 => x"5b5e0e4f",
  2213 => x"710e5d5c",
  2214 => x"87c8ff4b",
  2215 => x"48f4f0c2",
  2216 => x"497350c0",
  2217 => x"7087eae2",
  2218 => x"9cc24c49",
  2219 => x"cb49eecb",
  2220 => x"497087cc",
  2221 => x"f4f0c24d",
  2222 => x"c105bf97",
  2223 => x"66d087e2",
  2224 => x"fdf0c249",
  2225 => x"d60599bf",
  2226 => x"4966d487",
  2227 => x"bff5f0c2",
  2228 => x"87cb0599",
  2229 => x"f8e14973",
  2230 => x"02987087",
  2231 => x"c187c1c1",
  2232 => x"87c0fe4c",
  2233 => x"e1ca4975",
  2234 => x"02987087",
  2235 => x"f0c287c6",
  2236 => x"50c148f4",
  2237 => x"97f4f0c2",
  2238 => x"e3c005bf",
  2239 => x"fdf0c287",
  2240 => x"66d049bf",
  2241 => x"d6ff0599",
  2242 => x"f5f0c287",
  2243 => x"66d449bf",
  2244 => x"caff0599",
  2245 => x"e0497387",
  2246 => x"987087f7",
  2247 => x"87fffe05",
  2248 => x"dcfb4874",
  2249 => x"5b5e0e87",
  2250 => x"f40e5d5c",
  2251 => x"4c4dc086",
  2252 => x"c47ebfec",
  2253 => x"f1c248a6",
  2254 => x"c178bfc1",
  2255 => x"c71ec01e",
  2256 => x"87cdfd49",
  2257 => x"987086c8",
  2258 => x"ff87ce02",
  2259 => x"87ccfb49",
  2260 => x"ff49dac1",
  2261 => x"c187fadf",
  2262 => x"f4f0c24d",
  2263 => x"c302bf97",
  2264 => x"87c4d087",
  2265 => x"bff9f0c2",
  2266 => x"f6d5c24b",
  2267 => x"ebc005bf",
  2268 => x"49fdc387",
  2269 => x"87d9dfff",
  2270 => x"ff49fac3",
  2271 => x"7387d2df",
  2272 => x"99ffc349",
  2273 => x"49c01e71",
  2274 => x"7387cbfb",
  2275 => x"29b7c849",
  2276 => x"49c11e71",
  2277 => x"c887fffa",
  2278 => x"87c0c686",
  2279 => x"bffdf0c2",
  2280 => x"dd029b4b",
  2281 => x"f2d5c287",
  2282 => x"ddc749bf",
  2283 => x"05987087",
  2284 => x"4bc087c4",
  2285 => x"e0c287d2",
  2286 => x"87c2c749",
  2287 => x"58f6d5c2",
  2288 => x"d5c287c6",
  2289 => x"78c048f2",
  2290 => x"99c24973",
  2291 => x"c387ce05",
  2292 => x"ddff49eb",
  2293 => x"497087fb",
  2294 => x"c20299c2",
  2295 => x"734cfb87",
  2296 => x"0599c149",
  2297 => x"f4c387ce",
  2298 => x"e4ddff49",
  2299 => x"c2497087",
  2300 => x"87c20299",
  2301 => x"49734cfa",
  2302 => x"ce0599c8",
  2303 => x"49f5c387",
  2304 => x"87cdddff",
  2305 => x"99c24970",
  2306 => x"c287d502",
  2307 => x"02bfc5f1",
  2308 => x"c14887ca",
  2309 => x"c9f1c288",
  2310 => x"87c2c058",
  2311 => x"4dc14cff",
  2312 => x"99c44973",
  2313 => x"c387ce05",
  2314 => x"dcff49f2",
  2315 => x"497087e3",
  2316 => x"dc0299c2",
  2317 => x"c5f1c287",
  2318 => x"c7487ebf",
  2319 => x"c003a8b7",
  2320 => x"486e87cb",
  2321 => x"f1c280c1",
  2322 => x"c2c058c9",
  2323 => x"c14cfe87",
  2324 => x"49fdc34d",
  2325 => x"87f9dbff",
  2326 => x"99c24970",
  2327 => x"c287d502",
  2328 => x"02bfc5f1",
  2329 => x"c287c9c0",
  2330 => x"c048c5f1",
  2331 => x"87c2c078",
  2332 => x"4dc14cfd",
  2333 => x"ff49fac3",
  2334 => x"7087d6db",
  2335 => x"0299c249",
  2336 => x"c287d9c0",
  2337 => x"48bfc5f1",
  2338 => x"03a8b7c7",
  2339 => x"c287c9c0",
  2340 => x"c748c5f1",
  2341 => x"87c2c078",
  2342 => x"4dc14cfc",
  2343 => x"03acb7c0",
  2344 => x"c487d1c0",
  2345 => x"d8c14a66",
  2346 => x"c0026a82",
  2347 => x"4b6a87c6",
  2348 => x"0f734974",
  2349 => x"f0c31ec0",
  2350 => x"49dac11e",
  2351 => x"c887d2f7",
  2352 => x"02987086",
  2353 => x"c887e2c0",
  2354 => x"f1c248a6",
  2355 => x"c878bfc5",
  2356 => x"91cb4966",
  2357 => x"714866c4",
  2358 => x"6e7e7080",
  2359 => x"c8c002bf",
  2360 => x"4bbf6e87",
  2361 => x"734966c8",
  2362 => x"029d750f",
  2363 => x"c287c8c0",
  2364 => x"49bfc5f1",
  2365 => x"c287c0f3",
  2366 => x"02bffad5",
  2367 => x"4987ddc0",
  2368 => x"7087c7c2",
  2369 => x"d3c00298",
  2370 => x"c5f1c287",
  2371 => x"e6f249bf",
  2372 => x"f449c087",
  2373 => x"d5c287c6",
  2374 => x"78c048fa",
  2375 => x"e0f38ef4",
  2376 => x"5b5e0e87",
  2377 => x"1e0e5d5c",
  2378 => x"f1c24c71",
  2379 => x"c149bfc1",
  2380 => x"c14da1cd",
  2381 => x"7e6981d1",
  2382 => x"cf029c74",
  2383 => x"4ba5c487",
  2384 => x"f1c27b74",
  2385 => x"f249bfc1",
  2386 => x"7b6e87ff",
  2387 => x"c4059c74",
  2388 => x"c24bc087",
  2389 => x"734bc187",
  2390 => x"87c0f349",
  2391 => x"c70266d4",
  2392 => x"87da4987",
  2393 => x"87c24a70",
  2394 => x"d5c24ac0",
  2395 => x"f2265afe",
  2396 => x"000087cf",
  2397 => x"00000000",
  2398 => x"00000000",
  2399 => x"711e0000",
  2400 => x"bfc8ff4a",
  2401 => x"48a17249",
  2402 => x"ff1e4f26",
  2403 => x"fe89bfc8",
  2404 => x"c0c0c0c0",
  2405 => x"c401a9c0",
  2406 => x"c24ac087",
  2407 => x"724ac187",
  2408 => x"0e4f2648",
  2409 => x"5d5c5b5e",
  2410 => x"ff4b710e",
  2411 => x"66d04cd4",
  2412 => x"d678c048",
  2413 => x"d0d8ff49",
  2414 => x"7cffc387",
  2415 => x"ffc3496c",
  2416 => x"494d7199",
  2417 => x"c199f0c3",
  2418 => x"cb05a9e0",
  2419 => x"7cffc387",
  2420 => x"98c3486c",
  2421 => x"780866d0",
  2422 => x"6c7cffc3",
  2423 => x"31c8494a",
  2424 => x"6c7cffc3",
  2425 => x"72b2714a",
  2426 => x"c331c849",
  2427 => x"4a6c7cff",
  2428 => x"4972b271",
  2429 => x"ffc331c8",
  2430 => x"714a6c7c",
  2431 => x"48d0ffb2",
  2432 => x"7378e0c0",
  2433 => x"87c2029b",
  2434 => x"48757b72",
  2435 => x"4c264d26",
  2436 => x"4f264b26",
  2437 => x"0e4f261e",
  2438 => x"0e5c5b5e",
  2439 => x"1e7686f8",
  2440 => x"fd49a6c8",
  2441 => x"86c487fd",
  2442 => x"486e4b70",
  2443 => x"c203a8c2",
  2444 => x"4a7387f0",
  2445 => x"c19af0c3",
  2446 => x"c702aad0",
  2447 => x"aae0c187",
  2448 => x"87dec205",
  2449 => x"99c84973",
  2450 => x"ff87c302",
  2451 => x"4c7387c6",
  2452 => x"acc29cc3",
  2453 => x"87c2c105",
  2454 => x"c94966c4",
  2455 => x"c41e7131",
  2456 => x"92d44a66",
  2457 => x"49c9f1c2",
  2458 => x"cdfe8172",
  2459 => x"49d887f2",
  2460 => x"87d5d5ff",
  2461 => x"c21ec0c8",
  2462 => x"fd49e2df",
  2463 => x"ff87ede9",
  2464 => x"e0c048d0",
  2465 => x"e2dfc278",
  2466 => x"4a66cc1e",
  2467 => x"f1c292d4",
  2468 => x"817249c9",
  2469 => x"87f9cbfe",
  2470 => x"acc186cc",
  2471 => x"87c2c105",
  2472 => x"c94966c4",
  2473 => x"c41e7131",
  2474 => x"92d44a66",
  2475 => x"49c9f1c2",
  2476 => x"ccfe8172",
  2477 => x"dfc287ea",
  2478 => x"66c81ee2",
  2479 => x"c292d44a",
  2480 => x"7249c9f1",
  2481 => x"f9c9fe81",
  2482 => x"ff49d787",
  2483 => x"c887fad3",
  2484 => x"dfc21ec0",
  2485 => x"e7fd49e2",
  2486 => x"86cc87eb",
  2487 => x"c048d0ff",
  2488 => x"8ef878e0",
  2489 => x"0e87e7fc",
  2490 => x"5d5c5b5e",
  2491 => x"4d711e0e",
  2492 => x"d44cd4ff",
  2493 => x"c3487e66",
  2494 => x"c506a8b7",
  2495 => x"c148c087",
  2496 => x"497587e2",
  2497 => x"87fedafe",
  2498 => x"66c41e75",
  2499 => x"c293d44b",
  2500 => x"7383c9f1",
  2501 => x"d4c5fe49",
  2502 => x"6b83c887",
  2503 => x"48d0ff4b",
  2504 => x"dd78e1c8",
  2505 => x"c349737c",
  2506 => x"7c7199ff",
  2507 => x"b7c84973",
  2508 => x"99ffc329",
  2509 => x"49737c71",
  2510 => x"c329b7d0",
  2511 => x"7c7199ff",
  2512 => x"b7d84973",
  2513 => x"c07c7129",
  2514 => x"7c7c7c7c",
  2515 => x"7c7c7c7c",
  2516 => x"7c7c7c7c",
  2517 => x"c478e0c0",
  2518 => x"49dc1e66",
  2519 => x"87ced2ff",
  2520 => x"487386c8",
  2521 => x"87e4fa26",
  2522 => x"f6dec21e",
  2523 => x"b9c149bf",
  2524 => x"59fadec2",
  2525 => x"c348d4ff",
  2526 => x"d0ff78ff",
  2527 => x"78e1c848",
  2528 => x"c148d4ff",
  2529 => x"7131c478",
  2530 => x"48d0ff78",
  2531 => x"2678e0c0",
  2532 => x"dec21e4f",
  2533 => x"ecc21eea",
  2534 => x"c3fe49d8",
  2535 => x"86c487cf",
  2536 => x"c3029870",
  2537 => x"87c0ff87",
  2538 => x"35314f26",
  2539 => x"205a484b",
  2540 => x"46432020",
  2541 => x"00000047",
  2542 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
