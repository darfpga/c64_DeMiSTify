
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"7f",x"61",x"41",x"7f"),
     1 => (x"00",x"00",x"40",x"7e"),
     2 => (x"19",x"09",x"7f",x"7f"),
     3 => (x"00",x"00",x"66",x"7f"),
     4 => (x"59",x"4d",x"6f",x"26"),
     5 => (x"00",x"00",x"32",x"7b"),
     6 => (x"7f",x"7f",x"01",x"01"),
     7 => (x"00",x"00",x"01",x"01"),
     8 => (x"40",x"40",x"7f",x"3f"),
     9 => (x"00",x"00",x"3f",x"7f"),
    10 => (x"70",x"70",x"3f",x"0f"),
    11 => (x"7f",x"00",x"0f",x"3f"),
    12 => (x"30",x"18",x"30",x"7f"),
    13 => (x"41",x"00",x"7f",x"7f"),
    14 => (x"1c",x"1c",x"36",x"63"),
    15 => (x"01",x"41",x"63",x"36"),
    16 => (x"7c",x"7c",x"06",x"03"),
    17 => (x"61",x"01",x"03",x"06"),
    18 => (x"47",x"4d",x"59",x"71"),
    19 => (x"00",x"00",x"41",x"43"),
    20 => (x"41",x"7f",x"7f",x"00"),
    21 => (x"01",x"00",x"00",x"41"),
    22 => (x"18",x"0c",x"06",x"03"),
    23 => (x"00",x"40",x"60",x"30"),
    24 => (x"7f",x"41",x"41",x"00"),
    25 => (x"08",x"00",x"00",x"7f"),
    26 => (x"06",x"03",x"06",x"0c"),
    27 => (x"80",x"00",x"08",x"0c"),
    28 => (x"80",x"80",x"80",x"80"),
    29 => (x"00",x"00",x"80",x"80"),
    30 => (x"07",x"03",x"00",x"00"),
    31 => (x"00",x"00",x"00",x"04"),
    32 => (x"54",x"54",x"74",x"20"),
    33 => (x"00",x"00",x"78",x"7c"),
    34 => (x"44",x"44",x"7f",x"7f"),
    35 => (x"00",x"00",x"38",x"7c"),
    36 => (x"44",x"44",x"7c",x"38"),
    37 => (x"00",x"00",x"00",x"44"),
    38 => (x"44",x"44",x"7c",x"38"),
    39 => (x"00",x"00",x"7f",x"7f"),
    40 => (x"54",x"54",x"7c",x"38"),
    41 => (x"00",x"00",x"18",x"5c"),
    42 => (x"05",x"7f",x"7e",x"04"),
    43 => (x"00",x"00",x"00",x"05"),
    44 => (x"a4",x"a4",x"bc",x"18"),
    45 => (x"00",x"00",x"7c",x"fc"),
    46 => (x"04",x"04",x"7f",x"7f"),
    47 => (x"00",x"00",x"78",x"7c"),
    48 => (x"7d",x"3d",x"00",x"00"),
    49 => (x"00",x"00",x"00",x"40"),
    50 => (x"fd",x"80",x"80",x"80"),
    51 => (x"00",x"00",x"00",x"7d"),
    52 => (x"38",x"10",x"7f",x"7f"),
    53 => (x"00",x"00",x"44",x"6c"),
    54 => (x"7f",x"3f",x"00",x"00"),
    55 => (x"7c",x"00",x"00",x"40"),
    56 => (x"0c",x"18",x"0c",x"7c"),
    57 => (x"00",x"00",x"78",x"7c"),
    58 => (x"04",x"04",x"7c",x"7c"),
    59 => (x"00",x"00",x"78",x"7c"),
    60 => (x"44",x"44",x"7c",x"38"),
    61 => (x"00",x"00",x"38",x"7c"),
    62 => (x"24",x"24",x"fc",x"fc"),
    63 => (x"00",x"00",x"18",x"3c"),
    64 => (x"24",x"24",x"3c",x"18"),
    65 => (x"00",x"00",x"fc",x"fc"),
    66 => (x"04",x"04",x"7c",x"7c"),
    67 => (x"00",x"00",x"08",x"0c"),
    68 => (x"54",x"54",x"5c",x"48"),
    69 => (x"00",x"00",x"20",x"74"),
    70 => (x"44",x"7f",x"3f",x"04"),
    71 => (x"00",x"00",x"00",x"44"),
    72 => (x"40",x"40",x"7c",x"3c"),
    73 => (x"00",x"00",x"7c",x"7c"),
    74 => (x"60",x"60",x"3c",x"1c"),
    75 => (x"3c",x"00",x"1c",x"3c"),
    76 => (x"60",x"30",x"60",x"7c"),
    77 => (x"44",x"00",x"3c",x"7c"),
    78 => (x"38",x"10",x"38",x"6c"),
    79 => (x"00",x"00",x"44",x"6c"),
    80 => (x"60",x"e0",x"bc",x"1c"),
    81 => (x"00",x"00",x"1c",x"3c"),
    82 => (x"5c",x"74",x"64",x"44"),
    83 => (x"00",x"00",x"44",x"4c"),
    84 => (x"77",x"3e",x"08",x"08"),
    85 => (x"00",x"00",x"41",x"41"),
    86 => (x"7f",x"7f",x"00",x"00"),
    87 => (x"00",x"00",x"00",x"00"),
    88 => (x"3e",x"77",x"41",x"41"),
    89 => (x"02",x"00",x"08",x"08"),
    90 => (x"02",x"03",x"01",x"01"),
    91 => (x"7f",x"00",x"01",x"02"),
    92 => (x"7f",x"7f",x"7f",x"7f"),
    93 => (x"08",x"00",x"7f",x"7f"),
    94 => (x"3e",x"1c",x"1c",x"08"),
    95 => (x"7f",x"7f",x"7f",x"3e"),
    96 => (x"1c",x"3e",x"3e",x"7f"),
    97 => (x"00",x"08",x"08",x"1c"),
    98 => (x"7c",x"7c",x"18",x"10"),
    99 => (x"00",x"00",x"10",x"18"),
   100 => (x"7c",x"7c",x"30",x"10"),
   101 => (x"10",x"00",x"10",x"30"),
   102 => (x"78",x"60",x"60",x"30"),
   103 => (x"42",x"00",x"06",x"1e"),
   104 => (x"3c",x"18",x"3c",x"66"),
   105 => (x"78",x"00",x"42",x"66"),
   106 => (x"c6",x"c2",x"6a",x"38"),
   107 => (x"60",x"00",x"38",x"6c"),
   108 => (x"00",x"60",x"00",x"00"),
   109 => (x"0e",x"00",x"60",x"00"),
   110 => (x"5d",x"5c",x"5b",x"5e"),
   111 => (x"4c",x"71",x"1e",x"0e"),
   112 => (x"bf",x"c1",x"f1",x"c2"),
   113 => (x"c0",x"4b",x"c0",x"4d"),
   114 => (x"02",x"ab",x"74",x"1e"),
   115 => (x"a6",x"c4",x"87",x"c7"),
   116 => (x"c5",x"78",x"c0",x"48"),
   117 => (x"48",x"a6",x"c4",x"87"),
   118 => (x"66",x"c4",x"78",x"c1"),
   119 => (x"ee",x"49",x"73",x"1e"),
   120 => (x"86",x"c8",x"87",x"df"),
   121 => (x"ef",x"49",x"e0",x"c0"),
   122 => (x"a5",x"c4",x"87",x"ef"),
   123 => (x"f0",x"49",x"6a",x"4a"),
   124 => (x"c6",x"f1",x"87",x"f0"),
   125 => (x"c1",x"85",x"cb",x"87"),
   126 => (x"ab",x"b7",x"c8",x"83"),
   127 => (x"87",x"c7",x"ff",x"04"),
   128 => (x"26",x"4d",x"26",x"26"),
   129 => (x"26",x"4b",x"26",x"4c"),
   130 => (x"4a",x"71",x"1e",x"4f"),
   131 => (x"5a",x"c5",x"f1",x"c2"),
   132 => (x"48",x"c5",x"f1",x"c2"),
   133 => (x"fe",x"49",x"78",x"c7"),
   134 => (x"4f",x"26",x"87",x"dd"),
   135 => (x"71",x"1e",x"73",x"1e"),
   136 => (x"aa",x"b7",x"c0",x"4a"),
   137 => (x"c2",x"87",x"d3",x"03"),
   138 => (x"05",x"bf",x"f6",x"d5"),
   139 => (x"4b",x"c1",x"87",x"c4"),
   140 => (x"4b",x"c0",x"87",x"c2"),
   141 => (x"5b",x"fa",x"d5",x"c2"),
   142 => (x"d5",x"c2",x"87",x"c4"),
   143 => (x"d5",x"c2",x"5a",x"fa"),
   144 => (x"c1",x"4a",x"bf",x"f6"),
   145 => (x"a2",x"c0",x"c1",x"9a"),
   146 => (x"87",x"e8",x"ec",x"49"),
   147 => (x"d5",x"c2",x"48",x"fc"),
   148 => (x"fe",x"78",x"bf",x"f6"),
   149 => (x"71",x"1e",x"87",x"ef"),
   150 => (x"1e",x"66",x"c4",x"4a"),
   151 => (x"e2",x"e6",x"49",x"72"),
   152 => (x"4f",x"26",x"26",x"87"),
   153 => (x"f6",x"d5",x"c2",x"1e"),
   154 => (x"c4",x"e3",x"49",x"bf"),
   155 => (x"f9",x"f0",x"c2",x"87"),
   156 => (x"78",x"bf",x"e8",x"48"),
   157 => (x"48",x"f5",x"f0",x"c2"),
   158 => (x"c2",x"78",x"bf",x"ec"),
   159 => (x"4a",x"bf",x"f9",x"f0"),
   160 => (x"99",x"ff",x"c3",x"49"),
   161 => (x"72",x"2a",x"b7",x"c8"),
   162 => (x"c2",x"b0",x"71",x"48"),
   163 => (x"26",x"58",x"c1",x"f1"),
   164 => (x"5b",x"5e",x"0e",x"4f"),
   165 => (x"71",x"0e",x"5d",x"5c"),
   166 => (x"87",x"c8",x"ff",x"4b"),
   167 => (x"48",x"f4",x"f0",x"c2"),
   168 => (x"49",x"73",x"50",x"c0"),
   169 => (x"70",x"87",x"ea",x"e2"),
   170 => (x"9c",x"c2",x"4c",x"49"),
   171 => (x"cb",x"49",x"ee",x"cb"),
   172 => (x"49",x"70",x"87",x"cc"),
   173 => (x"f4",x"f0",x"c2",x"4d"),
   174 => (x"c1",x"05",x"bf",x"97"),
   175 => (x"66",x"d0",x"87",x"e2"),
   176 => (x"fd",x"f0",x"c2",x"49"),
   177 => (x"d6",x"05",x"99",x"bf"),
   178 => (x"49",x"66",x"d4",x"87"),
   179 => (x"bf",x"f5",x"f0",x"c2"),
   180 => (x"87",x"cb",x"05",x"99"),
   181 => (x"f8",x"e1",x"49",x"73"),
   182 => (x"02",x"98",x"70",x"87"),
   183 => (x"c1",x"87",x"c1",x"c1"),
   184 => (x"87",x"c0",x"fe",x"4c"),
   185 => (x"e1",x"ca",x"49",x"75"),
   186 => (x"02",x"98",x"70",x"87"),
   187 => (x"f0",x"c2",x"87",x"c6"),
   188 => (x"50",x"c1",x"48",x"f4"),
   189 => (x"97",x"f4",x"f0",x"c2"),
   190 => (x"e3",x"c0",x"05",x"bf"),
   191 => (x"fd",x"f0",x"c2",x"87"),
   192 => (x"66",x"d0",x"49",x"bf"),
   193 => (x"d6",x"ff",x"05",x"99"),
   194 => (x"f5",x"f0",x"c2",x"87"),
   195 => (x"66",x"d4",x"49",x"bf"),
   196 => (x"ca",x"ff",x"05",x"99"),
   197 => (x"e0",x"49",x"73",x"87"),
   198 => (x"98",x"70",x"87",x"f7"),
   199 => (x"87",x"ff",x"fe",x"05"),
   200 => (x"dc",x"fb",x"48",x"74"),
   201 => (x"5b",x"5e",x"0e",x"87"),
   202 => (x"f4",x"0e",x"5d",x"5c"),
   203 => (x"4c",x"4d",x"c0",x"86"),
   204 => (x"c4",x"7e",x"bf",x"ec"),
   205 => (x"f1",x"c2",x"48",x"a6"),
   206 => (x"c1",x"78",x"bf",x"c1"),
   207 => (x"c7",x"1e",x"c0",x"1e"),
   208 => (x"87",x"cd",x"fd",x"49"),
   209 => (x"98",x"70",x"86",x"c8"),
   210 => (x"ff",x"87",x"ce",x"02"),
   211 => (x"87",x"cc",x"fb",x"49"),
   212 => (x"ff",x"49",x"da",x"c1"),
   213 => (x"c1",x"87",x"fa",x"df"),
   214 => (x"f4",x"f0",x"c2",x"4d"),
   215 => (x"c3",x"02",x"bf",x"97"),
   216 => (x"87",x"c4",x"d0",x"87"),
   217 => (x"bf",x"f9",x"f0",x"c2"),
   218 => (x"f6",x"d5",x"c2",x"4b"),
   219 => (x"eb",x"c0",x"05",x"bf"),
   220 => (x"49",x"fd",x"c3",x"87"),
   221 => (x"87",x"d9",x"df",x"ff"),
   222 => (x"ff",x"49",x"fa",x"c3"),
   223 => (x"73",x"87",x"d2",x"df"),
   224 => (x"99",x"ff",x"c3",x"49"),
   225 => (x"49",x"c0",x"1e",x"71"),
   226 => (x"73",x"87",x"cb",x"fb"),
   227 => (x"29",x"b7",x"c8",x"49"),
   228 => (x"49",x"c1",x"1e",x"71"),
   229 => (x"c8",x"87",x"ff",x"fa"),
   230 => (x"87",x"c0",x"c6",x"86"),
   231 => (x"bf",x"fd",x"f0",x"c2"),
   232 => (x"dd",x"02",x"9b",x"4b"),
   233 => (x"f2",x"d5",x"c2",x"87"),
   234 => (x"dd",x"c7",x"49",x"bf"),
   235 => (x"05",x"98",x"70",x"87"),
   236 => (x"4b",x"c0",x"87",x"c4"),
   237 => (x"e0",x"c2",x"87",x"d2"),
   238 => (x"87",x"c2",x"c7",x"49"),
   239 => (x"58",x"f6",x"d5",x"c2"),
   240 => (x"d5",x"c2",x"87",x"c6"),
   241 => (x"78",x"c0",x"48",x"f2"),
   242 => (x"99",x"c2",x"49",x"73"),
   243 => (x"c3",x"87",x"ce",x"05"),
   244 => (x"dd",x"ff",x"49",x"eb"),
   245 => (x"49",x"70",x"87",x"fb"),
   246 => (x"c2",x"02",x"99",x"c2"),
   247 => (x"73",x"4c",x"fb",x"87"),
   248 => (x"05",x"99",x"c1",x"49"),
   249 => (x"f4",x"c3",x"87",x"ce"),
   250 => (x"e4",x"dd",x"ff",x"49"),
   251 => (x"c2",x"49",x"70",x"87"),
   252 => (x"87",x"c2",x"02",x"99"),
   253 => (x"49",x"73",x"4c",x"fa"),
   254 => (x"ce",x"05",x"99",x"c8"),
   255 => (x"49",x"f5",x"c3",x"87"),
   256 => (x"87",x"cd",x"dd",x"ff"),
   257 => (x"99",x"c2",x"49",x"70"),
   258 => (x"c2",x"87",x"d5",x"02"),
   259 => (x"02",x"bf",x"c5",x"f1"),
   260 => (x"c1",x"48",x"87",x"ca"),
   261 => (x"c9",x"f1",x"c2",x"88"),
   262 => (x"87",x"c2",x"c0",x"58"),
   263 => (x"4d",x"c1",x"4c",x"ff"),
   264 => (x"99",x"c4",x"49",x"73"),
   265 => (x"c3",x"87",x"ce",x"05"),
   266 => (x"dc",x"ff",x"49",x"f2"),
   267 => (x"49",x"70",x"87",x"e3"),
   268 => (x"dc",x"02",x"99",x"c2"),
   269 => (x"c5",x"f1",x"c2",x"87"),
   270 => (x"c7",x"48",x"7e",x"bf"),
   271 => (x"c0",x"03",x"a8",x"b7"),
   272 => (x"48",x"6e",x"87",x"cb"),
   273 => (x"f1",x"c2",x"80",x"c1"),
   274 => (x"c2",x"c0",x"58",x"c9"),
   275 => (x"c1",x"4c",x"fe",x"87"),
   276 => (x"49",x"fd",x"c3",x"4d"),
   277 => (x"87",x"f9",x"db",x"ff"),
   278 => (x"99",x"c2",x"49",x"70"),
   279 => (x"c2",x"87",x"d5",x"02"),
   280 => (x"02",x"bf",x"c5",x"f1"),
   281 => (x"c2",x"87",x"c9",x"c0"),
   282 => (x"c0",x"48",x"c5",x"f1"),
   283 => (x"87",x"c2",x"c0",x"78"),
   284 => (x"4d",x"c1",x"4c",x"fd"),
   285 => (x"ff",x"49",x"fa",x"c3"),
   286 => (x"70",x"87",x"d6",x"db"),
   287 => (x"02",x"99",x"c2",x"49"),
   288 => (x"c2",x"87",x"d9",x"c0"),
   289 => (x"48",x"bf",x"c5",x"f1"),
   290 => (x"03",x"a8",x"b7",x"c7"),
   291 => (x"c2",x"87",x"c9",x"c0"),
   292 => (x"c7",x"48",x"c5",x"f1"),
   293 => (x"87",x"c2",x"c0",x"78"),
   294 => (x"4d",x"c1",x"4c",x"fc"),
   295 => (x"03",x"ac",x"b7",x"c0"),
   296 => (x"c4",x"87",x"d1",x"c0"),
   297 => (x"d8",x"c1",x"4a",x"66"),
   298 => (x"c0",x"02",x"6a",x"82"),
   299 => (x"4b",x"6a",x"87",x"c6"),
   300 => (x"0f",x"73",x"49",x"74"),
   301 => (x"f0",x"c3",x"1e",x"c0"),
   302 => (x"49",x"da",x"c1",x"1e"),
   303 => (x"c8",x"87",x"d2",x"f7"),
   304 => (x"02",x"98",x"70",x"86"),
   305 => (x"c8",x"87",x"e2",x"c0"),
   306 => (x"f1",x"c2",x"48",x"a6"),
   307 => (x"c8",x"78",x"bf",x"c5"),
   308 => (x"91",x"cb",x"49",x"66"),
   309 => (x"71",x"48",x"66",x"c4"),
   310 => (x"6e",x"7e",x"70",x"80"),
   311 => (x"c8",x"c0",x"02",x"bf"),
   312 => (x"4b",x"bf",x"6e",x"87"),
   313 => (x"73",x"49",x"66",x"c8"),
   314 => (x"02",x"9d",x"75",x"0f"),
   315 => (x"c2",x"87",x"c8",x"c0"),
   316 => (x"49",x"bf",x"c5",x"f1"),
   317 => (x"c2",x"87",x"c0",x"f3"),
   318 => (x"02",x"bf",x"fa",x"d5"),
   319 => (x"49",x"87",x"dd",x"c0"),
   320 => (x"70",x"87",x"c7",x"c2"),
   321 => (x"d3",x"c0",x"02",x"98"),
   322 => (x"c5",x"f1",x"c2",x"87"),
   323 => (x"e6",x"f2",x"49",x"bf"),
   324 => (x"f4",x"49",x"c0",x"87"),
   325 => (x"d5",x"c2",x"87",x"c6"),
   326 => (x"78",x"c0",x"48",x"fa"),
   327 => (x"e0",x"f3",x"8e",x"f4"),
   328 => (x"5b",x"5e",x"0e",x"87"),
   329 => (x"1e",x"0e",x"5d",x"5c"),
   330 => (x"f1",x"c2",x"4c",x"71"),
   331 => (x"c1",x"49",x"bf",x"c1"),
   332 => (x"c1",x"4d",x"a1",x"cd"),
   333 => (x"7e",x"69",x"81",x"d1"),
   334 => (x"cf",x"02",x"9c",x"74"),
   335 => (x"4b",x"a5",x"c4",x"87"),
   336 => (x"f1",x"c2",x"7b",x"74"),
   337 => (x"f2",x"49",x"bf",x"c1"),
   338 => (x"7b",x"6e",x"87",x"ff"),
   339 => (x"c4",x"05",x"9c",x"74"),
   340 => (x"c2",x"4b",x"c0",x"87"),
   341 => (x"73",x"4b",x"c1",x"87"),
   342 => (x"87",x"c0",x"f3",x"49"),
   343 => (x"c7",x"02",x"66",x"d4"),
   344 => (x"87",x"da",x"49",x"87"),
   345 => (x"87",x"c2",x"4a",x"70"),
   346 => (x"d5",x"c2",x"4a",x"c0"),
   347 => (x"f2",x"26",x"5a",x"fe"),
   348 => (x"00",x"00",x"87",x"cf"),
   349 => (x"00",x"00",x"00",x"00"),
   350 => (x"00",x"00",x"00",x"00"),
   351 => (x"71",x"1e",x"00",x"00"),
   352 => (x"bf",x"c8",x"ff",x"4a"),
   353 => (x"48",x"a1",x"72",x"49"),
   354 => (x"ff",x"1e",x"4f",x"26"),
   355 => (x"fe",x"89",x"bf",x"c8"),
   356 => (x"c0",x"c0",x"c0",x"c0"),
   357 => (x"c4",x"01",x"a9",x"c0"),
   358 => (x"c2",x"4a",x"c0",x"87"),
   359 => (x"72",x"4a",x"c1",x"87"),
   360 => (x"0e",x"4f",x"26",x"48"),
   361 => (x"5d",x"5c",x"5b",x"5e"),
   362 => (x"ff",x"4b",x"71",x"0e"),
   363 => (x"66",x"d0",x"4c",x"d4"),
   364 => (x"d6",x"78",x"c0",x"48"),
   365 => (x"d0",x"d8",x"ff",x"49"),
   366 => (x"7c",x"ff",x"c3",x"87"),
   367 => (x"ff",x"c3",x"49",x"6c"),
   368 => (x"49",x"4d",x"71",x"99"),
   369 => (x"c1",x"99",x"f0",x"c3"),
   370 => (x"cb",x"05",x"a9",x"e0"),
   371 => (x"7c",x"ff",x"c3",x"87"),
   372 => (x"98",x"c3",x"48",x"6c"),
   373 => (x"78",x"08",x"66",x"d0"),
   374 => (x"6c",x"7c",x"ff",x"c3"),
   375 => (x"31",x"c8",x"49",x"4a"),
   376 => (x"6c",x"7c",x"ff",x"c3"),
   377 => (x"72",x"b2",x"71",x"4a"),
   378 => (x"c3",x"31",x"c8",x"49"),
   379 => (x"4a",x"6c",x"7c",x"ff"),
   380 => (x"49",x"72",x"b2",x"71"),
   381 => (x"ff",x"c3",x"31",x"c8"),
   382 => (x"71",x"4a",x"6c",x"7c"),
   383 => (x"48",x"d0",x"ff",x"b2"),
   384 => (x"73",x"78",x"e0",x"c0"),
   385 => (x"87",x"c2",x"02",x"9b"),
   386 => (x"48",x"75",x"7b",x"72"),
   387 => (x"4c",x"26",x"4d",x"26"),
   388 => (x"4f",x"26",x"4b",x"26"),
   389 => (x"0e",x"4f",x"26",x"1e"),
   390 => (x"0e",x"5c",x"5b",x"5e"),
   391 => (x"1e",x"76",x"86",x"f8"),
   392 => (x"fd",x"49",x"a6",x"c8"),
   393 => (x"86",x"c4",x"87",x"fd"),
   394 => (x"48",x"6e",x"4b",x"70"),
   395 => (x"c2",x"03",x"a8",x"c2"),
   396 => (x"4a",x"73",x"87",x"f0"),
   397 => (x"c1",x"9a",x"f0",x"c3"),
   398 => (x"c7",x"02",x"aa",x"d0"),
   399 => (x"aa",x"e0",x"c1",x"87"),
   400 => (x"87",x"de",x"c2",x"05"),
   401 => (x"99",x"c8",x"49",x"73"),
   402 => (x"ff",x"87",x"c3",x"02"),
   403 => (x"4c",x"73",x"87",x"c6"),
   404 => (x"ac",x"c2",x"9c",x"c3"),
   405 => (x"87",x"c2",x"c1",x"05"),
   406 => (x"c9",x"49",x"66",x"c4"),
   407 => (x"c4",x"1e",x"71",x"31"),
   408 => (x"92",x"d4",x"4a",x"66"),
   409 => (x"49",x"c9",x"f1",x"c2"),
   410 => (x"cd",x"fe",x"81",x"72"),
   411 => (x"49",x"d8",x"87",x"f2"),
   412 => (x"87",x"d5",x"d5",x"ff"),
   413 => (x"c2",x"1e",x"c0",x"c8"),
   414 => (x"fd",x"49",x"e2",x"df"),
   415 => (x"ff",x"87",x"ed",x"e9"),
   416 => (x"e0",x"c0",x"48",x"d0"),
   417 => (x"e2",x"df",x"c2",x"78"),
   418 => (x"4a",x"66",x"cc",x"1e"),
   419 => (x"f1",x"c2",x"92",x"d4"),
   420 => (x"81",x"72",x"49",x"c9"),
   421 => (x"87",x"f9",x"cb",x"fe"),
   422 => (x"ac",x"c1",x"86",x"cc"),
   423 => (x"87",x"c2",x"c1",x"05"),
   424 => (x"c9",x"49",x"66",x"c4"),
   425 => (x"c4",x"1e",x"71",x"31"),
   426 => (x"92",x"d4",x"4a",x"66"),
   427 => (x"49",x"c9",x"f1",x"c2"),
   428 => (x"cc",x"fe",x"81",x"72"),
   429 => (x"df",x"c2",x"87",x"ea"),
   430 => (x"66",x"c8",x"1e",x"e2"),
   431 => (x"c2",x"92",x"d4",x"4a"),
   432 => (x"72",x"49",x"c9",x"f1"),
   433 => (x"f9",x"c9",x"fe",x"81"),
   434 => (x"ff",x"49",x"d7",x"87"),
   435 => (x"c8",x"87",x"fa",x"d3"),
   436 => (x"df",x"c2",x"1e",x"c0"),
   437 => (x"e7",x"fd",x"49",x"e2"),
   438 => (x"86",x"cc",x"87",x"eb"),
   439 => (x"c0",x"48",x"d0",x"ff"),
   440 => (x"8e",x"f8",x"78",x"e0"),
   441 => (x"0e",x"87",x"e7",x"fc"),
   442 => (x"5d",x"5c",x"5b",x"5e"),
   443 => (x"4d",x"71",x"1e",x"0e"),
   444 => (x"d4",x"4c",x"d4",x"ff"),
   445 => (x"c3",x"48",x"7e",x"66"),
   446 => (x"c5",x"06",x"a8",x"b7"),
   447 => (x"c1",x"48",x"c0",x"87"),
   448 => (x"49",x"75",x"87",x"e2"),
   449 => (x"87",x"fe",x"da",x"fe"),
   450 => (x"66",x"c4",x"1e",x"75"),
   451 => (x"c2",x"93",x"d4",x"4b"),
   452 => (x"73",x"83",x"c9",x"f1"),
   453 => (x"d4",x"c5",x"fe",x"49"),
   454 => (x"6b",x"83",x"c8",x"87"),
   455 => (x"48",x"d0",x"ff",x"4b"),
   456 => (x"dd",x"78",x"e1",x"c8"),
   457 => (x"c3",x"49",x"73",x"7c"),
   458 => (x"7c",x"71",x"99",x"ff"),
   459 => (x"b7",x"c8",x"49",x"73"),
   460 => (x"99",x"ff",x"c3",x"29"),
   461 => (x"49",x"73",x"7c",x"71"),
   462 => (x"c3",x"29",x"b7",x"d0"),
   463 => (x"7c",x"71",x"99",x"ff"),
   464 => (x"b7",x"d8",x"49",x"73"),
   465 => (x"c0",x"7c",x"71",x"29"),
   466 => (x"7c",x"7c",x"7c",x"7c"),
   467 => (x"7c",x"7c",x"7c",x"7c"),
   468 => (x"7c",x"7c",x"7c",x"7c"),
   469 => (x"c4",x"78",x"e0",x"c0"),
   470 => (x"49",x"dc",x"1e",x"66"),
   471 => (x"87",x"ce",x"d2",x"ff"),
   472 => (x"48",x"73",x"86",x"c8"),
   473 => (x"87",x"e4",x"fa",x"26"),
   474 => (x"f6",x"de",x"c2",x"1e"),
   475 => (x"b9",x"c1",x"49",x"bf"),
   476 => (x"59",x"fa",x"de",x"c2"),
   477 => (x"c3",x"48",x"d4",x"ff"),
   478 => (x"d0",x"ff",x"78",x"ff"),
   479 => (x"78",x"e1",x"c8",x"48"),
   480 => (x"c1",x"48",x"d4",x"ff"),
   481 => (x"71",x"31",x"c4",x"78"),
   482 => (x"48",x"d0",x"ff",x"78"),
   483 => (x"26",x"78",x"e0",x"c0"),
   484 => (x"de",x"c2",x"1e",x"4f"),
   485 => (x"ec",x"c2",x"1e",x"ea"),
   486 => (x"c3",x"fe",x"49",x"d8"),
   487 => (x"86",x"c4",x"87",x"cf"),
   488 => (x"c3",x"02",x"98",x"70"),
   489 => (x"87",x"c0",x"ff",x"87"),
   490 => (x"35",x"31",x"4f",x"26"),
   491 => (x"20",x"5a",x"48",x"4b"),
   492 => (x"46",x"43",x"20",x"20"),
   493 => (x"00",x"00",x"00",x"47"),
   494 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

