library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"dce0c287",
    12 => x"86c0c84e",
    13 => x"49dce0c2",
    14 => x"48d0cec2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087d2dc",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"c44a711e",
    47 => x"c1484966",
    48 => x"58a6c888",
    49 => x"d6029971",
    50 => x"48d4ff87",
    51 => x"6878ffc3",
    52 => x"4966c452",
    53 => x"c888c148",
    54 => x"997158a6",
    55 => x"2687ea05",
    56 => x"1e731e4f",
    57 => x"c34bd4ff",
    58 => x"4a6b7bff",
    59 => x"6b7bffc3",
    60 => x"7232c849",
    61 => x"7bffc3b1",
    62 => x"31c84a6b",
    63 => x"ffc3b271",
    64 => x"c8496b7b",
    65 => x"71b17232",
    66 => x"2687c448",
    67 => x"264c264d",
    68 => x"0e4f264b",
    69 => x"5d5c5b5e",
    70 => x"ff4a710e",
    71 => x"49724cd4",
    72 => x"7199ffc3",
    73 => x"d0cec27c",
    74 => x"87c805bf",
    75 => x"c94866d0",
    76 => x"58a6d430",
    77 => x"d84966d0",
    78 => x"99ffc329",
    79 => x"66d07c71",
    80 => x"c329d049",
    81 => x"7c7199ff",
    82 => x"c84966d0",
    83 => x"99ffc329",
    84 => x"66d07c71",
    85 => x"99ffc349",
    86 => x"49727c71",
    87 => x"ffc329d0",
    88 => x"6c7c7199",
    89 => x"fff0c94b",
    90 => x"abffc34d",
    91 => x"c387d005",
    92 => x"4b6c7cff",
    93 => x"c6028dc1",
    94 => x"abffc387",
    95 => x"7387f002",
    96 => x"87c7fe48",
    97 => x"ff49c01e",
    98 => x"ffc348d4",
    99 => x"c381c178",
   100 => x"04a9b7c8",
   101 => x"4f2687f1",
   102 => x"e71e731e",
   103 => x"dff8c487",
   104 => x"c01ec04b",
   105 => x"f7c1f0ff",
   106 => x"87e7fd49",
   107 => x"a8c186c4",
   108 => x"87eac005",
   109 => x"c348d4ff",
   110 => x"c0c178ff",
   111 => x"c0c0c0c0",
   112 => x"f0e1c01e",
   113 => x"fd49e9c1",
   114 => x"86c487c9",
   115 => x"ca059870",
   116 => x"48d4ff87",
   117 => x"c178ffc3",
   118 => x"fe87cb48",
   119 => x"8bc187e6",
   120 => x"87fdfe05",
   121 => x"e6fc48c0",
   122 => x"1e731e87",
   123 => x"c348d4ff",
   124 => x"4bd378ff",
   125 => x"ffc01ec0",
   126 => x"49c1c1f0",
   127 => x"c487d4fc",
   128 => x"05987086",
   129 => x"d4ff87ca",
   130 => x"78ffc348",
   131 => x"87cb48c1",
   132 => x"c187f1fd",
   133 => x"dbff058b",
   134 => x"fb48c087",
   135 => x"5e0e87f1",
   136 => x"ff0e5c5b",
   137 => x"dbfd4cd4",
   138 => x"1eeac687",
   139 => x"c1f0e1c0",
   140 => x"defb49c8",
   141 => x"c186c487",
   142 => x"87c802a8",
   143 => x"c087eafe",
   144 => x"87e2c148",
   145 => x"7087dafa",
   146 => x"ffffcf49",
   147 => x"a9eac699",
   148 => x"fe87c802",
   149 => x"48c087d3",
   150 => x"c387cbc1",
   151 => x"f1c07cff",
   152 => x"87f4fc4b",
   153 => x"c0029870",
   154 => x"1ec087eb",
   155 => x"c1f0ffc0",
   156 => x"defa49fa",
   157 => x"7086c487",
   158 => x"87d90598",
   159 => x"6c7cffc3",
   160 => x"7cffc349",
   161 => x"c17c7c7c",
   162 => x"c40299c0",
   163 => x"d548c187",
   164 => x"d148c087",
   165 => x"05abc287",
   166 => x"48c087c4",
   167 => x"8bc187c8",
   168 => x"87fdfe05",
   169 => x"e4f948c0",
   170 => x"1e731e87",
   171 => x"48d0cec2",
   172 => x"4bc778c1",
   173 => x"c248d0ff",
   174 => x"87c8fb78",
   175 => x"c348d0ff",
   176 => x"c01ec078",
   177 => x"c0c1d0e5",
   178 => x"87c7f949",
   179 => x"a8c186c4",
   180 => x"4b87c105",
   181 => x"c505abc2",
   182 => x"c048c087",
   183 => x"8bc187f9",
   184 => x"87d0ff05",
   185 => x"c287f7fc",
   186 => x"7058d4ce",
   187 => x"87cd0598",
   188 => x"ffc01ec1",
   189 => x"49d0c1f0",
   190 => x"c487d8f8",
   191 => x"48d4ff86",
   192 => x"c278ffc3",
   193 => x"cec287fc",
   194 => x"d0ff58d8",
   195 => x"ff78c248",
   196 => x"ffc348d4",
   197 => x"f748c178",
   198 => x"5e0e87f5",
   199 => x"0e5d5c5b",
   200 => x"4cc04b71",
   201 => x"dfcdeec5",
   202 => x"48d4ff4a",
   203 => x"6878ffc3",
   204 => x"a9fec349",
   205 => x"87fdc005",
   206 => x"9b734d70",
   207 => x"d087cc02",
   208 => x"49731e66",
   209 => x"c487f1f5",
   210 => x"ff87d686",
   211 => x"d1c448d0",
   212 => x"7dffc378",
   213 => x"c14866d0",
   214 => x"58a6d488",
   215 => x"f0059870",
   216 => x"48d4ff87",
   217 => x"7878ffc3",
   218 => x"c5059b73",
   219 => x"48d0ff87",
   220 => x"4ac178d0",
   221 => x"058ac14c",
   222 => x"7487eefe",
   223 => x"87cbf648",
   224 => x"711e731e",
   225 => x"ff4bc04a",
   226 => x"ffc348d4",
   227 => x"48d0ff78",
   228 => x"ff78c3c4",
   229 => x"ffc348d4",
   230 => x"c01e7278",
   231 => x"d1c1f0ff",
   232 => x"87eff549",
   233 => x"987086c4",
   234 => x"c887d205",
   235 => x"66cc1ec0",
   236 => x"87e6fd49",
   237 => x"4b7086c4",
   238 => x"c248d0ff",
   239 => x"f5487378",
   240 => x"5e0e87cd",
   241 => x"0e5d5c5b",
   242 => x"ffc01ec0",
   243 => x"49c9c1f0",
   244 => x"d287c0f5",
   245 => x"d8cec21e",
   246 => x"87fefc49",
   247 => x"4cc086c8",
   248 => x"b7d284c1",
   249 => x"87f804ac",
   250 => x"97d8cec2",
   251 => x"c0c349bf",
   252 => x"a9c0c199",
   253 => x"87e7c005",
   254 => x"97dfcec2",
   255 => x"31d049bf",
   256 => x"97e0cec2",
   257 => x"32c84abf",
   258 => x"cec2b172",
   259 => x"4abf97e1",
   260 => x"cf4c71b1",
   261 => x"9cffffff",
   262 => x"34ca84c1",
   263 => x"c287e7c1",
   264 => x"bf97e1ce",
   265 => x"c631c149",
   266 => x"e2cec299",
   267 => x"c74abf97",
   268 => x"b1722ab7",
   269 => x"97ddcec2",
   270 => x"cf4d4abf",
   271 => x"decec29d",
   272 => x"c34abf97",
   273 => x"c232ca9a",
   274 => x"bf97dfce",
   275 => x"7333c24b",
   276 => x"e0cec2b2",
   277 => x"c34bbf97",
   278 => x"b7c69bc0",
   279 => x"c2b2732b",
   280 => x"7148c181",
   281 => x"c1497030",
   282 => x"70307548",
   283 => x"c14c724d",
   284 => x"c8947184",
   285 => x"06adb7c0",
   286 => x"34c187cc",
   287 => x"c0c82db7",
   288 => x"ff01adb7",
   289 => x"487487f4",
   290 => x"0e87c0f2",
   291 => x"5d5c5b5e",
   292 => x"c286f80e",
   293 => x"c048fed6",
   294 => x"f6cec278",
   295 => x"fb49c01e",
   296 => x"86c487de",
   297 => x"c5059870",
   298 => x"c948c087",
   299 => x"4dc087ce",
   300 => x"edc07ec1",
   301 => x"c249bff3",
   302 => x"714aeccf",
   303 => x"e9ee4bc8",
   304 => x"05987087",
   305 => x"7ec087c2",
   306 => x"bfefedc0",
   307 => x"c8d0c249",
   308 => x"4bc8714a",
   309 => x"7087d3ee",
   310 => x"87c20598",
   311 => x"026e7ec0",
   312 => x"c287fdc0",
   313 => x"4dbffcd5",
   314 => x"9ff4d6c2",
   315 => x"c5487ebf",
   316 => x"05a8ead6",
   317 => x"d5c287c7",
   318 => x"ce4dbffc",
   319 => x"ca486e87",
   320 => x"02a8d5e9",
   321 => x"48c087c5",
   322 => x"c287f1c7",
   323 => x"751ef6ce",
   324 => x"87ecf949",
   325 => x"987086c4",
   326 => x"c087c505",
   327 => x"87dcc748",
   328 => x"bfefedc0",
   329 => x"c8d0c249",
   330 => x"4bc8714a",
   331 => x"7087fbec",
   332 => x"87c80598",
   333 => x"48fed6c2",
   334 => x"87da78c1",
   335 => x"bff3edc0",
   336 => x"eccfc249",
   337 => x"4bc8714a",
   338 => x"7087dfec",
   339 => x"c5c00298",
   340 => x"c648c087",
   341 => x"d6c287e6",
   342 => x"49bf97f4",
   343 => x"05a9d5c1",
   344 => x"c287cdc0",
   345 => x"bf97f5d6",
   346 => x"a9eac249",
   347 => x"87c5c002",
   348 => x"c7c648c0",
   349 => x"f6cec287",
   350 => x"487ebf97",
   351 => x"02a8e9c3",
   352 => x"6e87cec0",
   353 => x"a8ebc348",
   354 => x"87c5c002",
   355 => x"ebc548c0",
   356 => x"c1cfc287",
   357 => x"9949bf97",
   358 => x"87ccc005",
   359 => x"97c2cfc2",
   360 => x"a9c249bf",
   361 => x"87c5c002",
   362 => x"cfc548c0",
   363 => x"c3cfc287",
   364 => x"c248bf97",
   365 => x"7058fad6",
   366 => x"88c1484c",
   367 => x"58fed6c2",
   368 => x"97c4cfc2",
   369 => x"817549bf",
   370 => x"97c5cfc2",
   371 => x"32c84abf",
   372 => x"c27ea172",
   373 => x"6e48cbdb",
   374 => x"c6cfc278",
   375 => x"c848bf97",
   376 => x"d6c258a6",
   377 => x"c202bffe",
   378 => x"edc087d4",
   379 => x"c249bfef",
   380 => x"714ac8d0",
   381 => x"f1e94bc8",
   382 => x"02987087",
   383 => x"c087c5c0",
   384 => x"87f8c348",
   385 => x"bff6d6c2",
   386 => x"dfdbc24c",
   387 => x"dbcfc25c",
   388 => x"c849bf97",
   389 => x"dacfc231",
   390 => x"a14abf97",
   391 => x"dccfc249",
   392 => x"d04abf97",
   393 => x"49a17232",
   394 => x"97ddcfc2",
   395 => x"32d84abf",
   396 => x"c449a172",
   397 => x"dbc29166",
   398 => x"c281bfcb",
   399 => x"c259d3db",
   400 => x"bf97e3cf",
   401 => x"c232c84a",
   402 => x"bf97e2cf",
   403 => x"c24aa24b",
   404 => x"bf97e4cf",
   405 => x"7333d04b",
   406 => x"cfc24aa2",
   407 => x"4bbf97e5",
   408 => x"33d89bcf",
   409 => x"c24aa273",
   410 => x"c25ad7db",
   411 => x"4abfd3db",
   412 => x"92748ac2",
   413 => x"48d7dbc2",
   414 => x"c178a172",
   415 => x"cfc287ca",
   416 => x"49bf97c8",
   417 => x"cfc231c8",
   418 => x"4abf97c7",
   419 => x"d7c249a1",
   420 => x"d7c259c6",
   421 => x"c549bfc2",
   422 => x"81ffc731",
   423 => x"dbc229c9",
   424 => x"cfc259df",
   425 => x"4abf97cd",
   426 => x"cfc232c8",
   427 => x"4bbf97cc",
   428 => x"66c44aa2",
   429 => x"c2826e92",
   430 => x"c25adbdb",
   431 => x"c048d3db",
   432 => x"cfdbc278",
   433 => x"78a17248",
   434 => x"48dfdbc2",
   435 => x"bfd3dbc2",
   436 => x"e3dbc278",
   437 => x"d7dbc248",
   438 => x"d6c278bf",
   439 => x"c002bffe",
   440 => x"487487c9",
   441 => x"7e7030c4",
   442 => x"c287c9c0",
   443 => x"48bfdbdb",
   444 => x"7e7030c4",
   445 => x"48c2d7c2",
   446 => x"48c1786e",
   447 => x"4d268ef8",
   448 => x"4b264c26",
   449 => x"5e0e4f26",
   450 => x"0e5d5c5b",
   451 => x"d6c24a71",
   452 => x"cb02bffe",
   453 => x"c74b7287",
   454 => x"c14c722b",
   455 => x"87c99cff",
   456 => x"2bc84b72",
   457 => x"ffc34c72",
   458 => x"cbdbc29c",
   459 => x"edc083bf",
   460 => x"02abbfeb",
   461 => x"edc087d9",
   462 => x"cec25bef",
   463 => x"49731ef6",
   464 => x"c487fdf0",
   465 => x"05987086",
   466 => x"48c087c5",
   467 => x"c287e6c0",
   468 => x"02bffed6",
   469 => x"497487d2",
   470 => x"cec291c4",
   471 => x"4d6981f6",
   472 => x"ffffffcf",
   473 => x"87cb9dff",
   474 => x"91c24974",
   475 => x"81f6cec2",
   476 => x"754d699f",
   477 => x"87c6fe48",
   478 => x"5c5b5e0e",
   479 => x"86f80e5d",
   480 => x"059c4c71",
   481 => x"48c087c5",
   482 => x"c887c1c3",
   483 => x"486e7ea4",
   484 => x"66d878c0",
   485 => x"d887c702",
   486 => x"05bf9766",
   487 => x"48c087c5",
   488 => x"c087e9c2",
   489 => x"c749c11e",
   490 => x"86c487e6",
   491 => x"029d4d70",
   492 => x"c287c2c1",
   493 => x"d84ac6d7",
   494 => x"d2e24966",
   495 => x"02987087",
   496 => x"7587f2c0",
   497 => x"4966d84a",
   498 => x"f7e24bcb",
   499 => x"02987087",
   500 => x"c087e2c0",
   501 => x"029d751e",
   502 => x"a6c887c7",
   503 => x"c578c048",
   504 => x"48a6c887",
   505 => x"66c878c1",
   506 => x"87e4c649",
   507 => x"4d7086c4",
   508 => x"fefe059d",
   509 => x"029d7587",
   510 => x"dc87cfc1",
   511 => x"486e49a5",
   512 => x"a5da7869",
   513 => x"48a6c449",
   514 => x"9f78a4c4",
   515 => x"66c44869",
   516 => x"d6c27808",
   517 => x"d202bffe",
   518 => x"49a5d487",
   519 => x"c049699f",
   520 => x"7199ffff",
   521 => x"7030d048",
   522 => x"c087c27e",
   523 => x"48496e7e",
   524 => x"80bf66c4",
   525 => x"780866c4",
   526 => x"a4cc7cc0",
   527 => x"bf66c449",
   528 => x"49a4d079",
   529 => x"48c179c0",
   530 => x"48c087c2",
   531 => x"edfa8ef8",
   532 => x"5b5e0e87",
   533 => x"710e5d5c",
   534 => x"c1029c4c",
   535 => x"a4c887ca",
   536 => x"c1026949",
   537 => x"66d087c2",
   538 => x"82496c4a",
   539 => x"d05aa6d4",
   540 => x"c2b94d66",
   541 => x"4abffad6",
   542 => x"9972baff",
   543 => x"c0029971",
   544 => x"a4c487e4",
   545 => x"f9496b4b",
   546 => x"7b7087fc",
   547 => x"bff6d6c2",
   548 => x"71816c49",
   549 => x"c2b9757c",
   550 => x"4abffad6",
   551 => x"9972baff",
   552 => x"ff059971",
   553 => x"7c7587dc",
   554 => x"1e87d3f9",
   555 => x"4b711e73",
   556 => x"87c7029b",
   557 => x"6949a3c8",
   558 => x"c087c505",
   559 => x"87f7c048",
   560 => x"bfcfdbc2",
   561 => x"49a3c44a",
   562 => x"89c24969",
   563 => x"bff6d6c2",
   564 => x"4aa27191",
   565 => x"bffad6c2",
   566 => x"71996b49",
   567 => x"edc04aa2",
   568 => x"66c85aef",
   569 => x"ea49721e",
   570 => x"86c487d6",
   571 => x"c4059870",
   572 => x"c248c087",
   573 => x"f848c187",
   574 => x"731e87c8",
   575 => x"9b4b711e",
   576 => x"87e4c002",
   577 => x"5be3dbc2",
   578 => x"8ac24a73",
   579 => x"bff6d6c2",
   580 => x"dbc29249",
   581 => x"7248bfcf",
   582 => x"e7dbc280",
   583 => x"c4487158",
   584 => x"c6d7c230",
   585 => x"87edc058",
   586 => x"48dfdbc2",
   587 => x"bfd3dbc2",
   588 => x"e3dbc278",
   589 => x"d7dbc248",
   590 => x"d6c278bf",
   591 => x"c902bffe",
   592 => x"f6d6c287",
   593 => x"31c449bf",
   594 => x"dbc287c7",
   595 => x"c449bfdb",
   596 => x"c6d7c231",
   597 => x"87eaf659",
   598 => x"5c5b5e0e",
   599 => x"c04a710e",
   600 => x"029a724b",
   601 => x"da87e1c0",
   602 => x"699f49a2",
   603 => x"fed6c24b",
   604 => x"87cf02bf",
   605 => x"9f49a2d4",
   606 => x"c04c4969",
   607 => x"d09cffff",
   608 => x"c087c234",
   609 => x"b349744c",
   610 => x"edfd4973",
   611 => x"87f0f587",
   612 => x"5c5b5e0e",
   613 => x"86f40e5d",
   614 => x"7ec04a71",
   615 => x"d8029a72",
   616 => x"f2cec287",
   617 => x"c278c048",
   618 => x"c248eace",
   619 => x"78bfe3db",
   620 => x"48eecec2",
   621 => x"bfdfdbc2",
   622 => x"d3d7c278",
   623 => x"c250c048",
   624 => x"49bfc2d7",
   625 => x"bff2cec2",
   626 => x"03aa714a",
   627 => x"7287c9c4",
   628 => x"0599cf49",
   629 => x"c087e9c0",
   630 => x"c248ebed",
   631 => x"78bfeace",
   632 => x"1ef6cec2",
   633 => x"bfeacec2",
   634 => x"eacec249",
   635 => x"78a1c148",
   636 => x"87cce671",
   637 => x"edc086c4",
   638 => x"cec248e7",
   639 => x"87cc78f6",
   640 => x"bfe7edc0",
   641 => x"80e0c048",
   642 => x"58ebedc0",
   643 => x"bff2cec2",
   644 => x"c280c148",
   645 => x"2758f6ce",
   646 => x"00000b67",
   647 => x"4dbf97bf",
   648 => x"e3c2029d",
   649 => x"ade5c387",
   650 => x"87dcc202",
   651 => x"bfe7edc0",
   652 => x"49a3cb4b",
   653 => x"accf4c11",
   654 => x"87d2c105",
   655 => x"99df4975",
   656 => x"91cd89c1",
   657 => x"81c6d7c2",
   658 => x"124aa3c1",
   659 => x"4aa3c351",
   660 => x"a3c55112",
   661 => x"c751124a",
   662 => x"51124aa3",
   663 => x"124aa3c9",
   664 => x"4aa3ce51",
   665 => x"a3d05112",
   666 => x"d251124a",
   667 => x"51124aa3",
   668 => x"124aa3d4",
   669 => x"4aa3d651",
   670 => x"a3d85112",
   671 => x"dc51124a",
   672 => x"51124aa3",
   673 => x"124aa3de",
   674 => x"c07ec151",
   675 => x"497487fa",
   676 => x"c00599c8",
   677 => x"497487eb",
   678 => x"d10599d0",
   679 => x"0266dc87",
   680 => x"7387cbc0",
   681 => x"0f66dc49",
   682 => x"c0029870",
   683 => x"056e87d3",
   684 => x"c287c6c0",
   685 => x"c048c6d7",
   686 => x"e7edc050",
   687 => x"e1c248bf",
   688 => x"d3d7c287",
   689 => x"7e50c048",
   690 => x"bfc2d7c2",
   691 => x"f2cec249",
   692 => x"aa714abf",
   693 => x"87f7fb04",
   694 => x"bfe3dbc2",
   695 => x"87c8c005",
   696 => x"bffed6c2",
   697 => x"87f8c102",
   698 => x"bfeecec2",
   699 => x"87d6f049",
   700 => x"cec24970",
   701 => x"a6c459f2",
   702 => x"eecec248",
   703 => x"d6c278bf",
   704 => x"c002bffe",
   705 => x"66c487d8",
   706 => x"ffffcf49",
   707 => x"a999f8ff",
   708 => x"87c5c002",
   709 => x"e1c04cc0",
   710 => x"c04cc187",
   711 => x"66c487dc",
   712 => x"f8ffcf49",
   713 => x"c002a999",
   714 => x"a6c887c8",
   715 => x"c078c048",
   716 => x"a6c887c5",
   717 => x"c878c148",
   718 => x"9c744c66",
   719 => x"87e0c005",
   720 => x"c24966c4",
   721 => x"f6d6c289",
   722 => x"c2914abf",
   723 => x"4abfcfdb",
   724 => x"48eacec2",
   725 => x"c278a172",
   726 => x"c048f2ce",
   727 => x"87dff978",
   728 => x"8ef448c0",
   729 => x"0087d7ee",
   730 => x"ff000000",
   731 => x"77ffffff",
   732 => x"8000000b",
   733 => x"4600000b",
   734 => x"32335441",
   735 => x"00202020",
   736 => x"31544146",
   737 => x"20202036",
   738 => x"d4ff1e00",
   739 => x"78ffc348",
   740 => x"4f264868",
   741 => x"48d4ff1e",
   742 => x"ff78ffc3",
   743 => x"e1c048d0",
   744 => x"48d4ff78",
   745 => x"dbc278d4",
   746 => x"d4ff48e7",
   747 => x"4f2650bf",
   748 => x"48d0ff1e",
   749 => x"2678e0c0",
   750 => x"ccff1e4f",
   751 => x"99497087",
   752 => x"c087c602",
   753 => x"f105a9fb",
   754 => x"26487187",
   755 => x"5b5e0e4f",
   756 => x"4b710e5c",
   757 => x"f0fe4cc0",
   758 => x"99497087",
   759 => x"87f9c002",
   760 => x"02a9ecc0",
   761 => x"c087f2c0",
   762 => x"c002a9fb",
   763 => x"66cc87eb",
   764 => x"c703acb7",
   765 => x"0266d087",
   766 => x"537187c2",
   767 => x"c2029971",
   768 => x"fe84c187",
   769 => x"497087c3",
   770 => x"87cd0299",
   771 => x"02a9ecc0",
   772 => x"fbc087c7",
   773 => x"d5ff05a9",
   774 => x"0266d087",
   775 => x"97c087c3",
   776 => x"a9ecc07b",
   777 => x"7487c405",
   778 => x"7487c54a",
   779 => x"8a0ac04a",
   780 => x"87c24872",
   781 => x"4c264d26",
   782 => x"4f264b26",
   783 => x"87c9fd1e",
   784 => x"c04a4970",
   785 => x"c904aaf0",
   786 => x"aaf9c087",
   787 => x"c087c301",
   788 => x"c1c18af0",
   789 => x"87c904aa",
   790 => x"01aadac1",
   791 => x"f7c087c3",
   792 => x"2648728a",
   793 => x"5b5e0e4f",
   794 => x"4a710e5c",
   795 => x"724cd4ff",
   796 => x"87e9c049",
   797 => x"029b4b70",
   798 => x"8bc187c2",
   799 => x"c548d0ff",
   800 => x"7cd5c178",
   801 => x"31c64973",
   802 => x"97f3ddc1",
   803 => x"71484abf",
   804 => x"ff7c70b0",
   805 => x"78c448d0",
   806 => x"d9fe4873",
   807 => x"5b5e0e87",
   808 => x"f80e5d5c",
   809 => x"c04c7186",
   810 => x"87e8fb7e",
   811 => x"f5c04bc0",
   812 => x"49bf97ca",
   813 => x"cf04a9c0",
   814 => x"87fdfb87",
   815 => x"f5c083c1",
   816 => x"49bf97ca",
   817 => x"87f106ab",
   818 => x"97caf5c0",
   819 => x"87cf02bf",
   820 => x"7087f6fa",
   821 => x"c6029949",
   822 => x"a9ecc087",
   823 => x"c087f105",
   824 => x"87e5fa4b",
   825 => x"e0fa4d70",
   826 => x"58a6c887",
   827 => x"7087dafa",
   828 => x"c883c14a",
   829 => x"699749a4",
   830 => x"c702ad49",
   831 => x"adffc087",
   832 => x"87e7c005",
   833 => x"9749a4c9",
   834 => x"66c44969",
   835 => x"87c702a9",
   836 => x"a8ffc048",
   837 => x"ca87d405",
   838 => x"699749a4",
   839 => x"c602aa49",
   840 => x"aaffc087",
   841 => x"c187c405",
   842 => x"c087d07e",
   843 => x"c602adec",
   844 => x"adfbc087",
   845 => x"c087c405",
   846 => x"6e7ec14b",
   847 => x"87e1fe02",
   848 => x"7387edf9",
   849 => x"fb8ef848",
   850 => x"0e0087ea",
   851 => x"5d5c5b5e",
   852 => x"7186f80e",
   853 => x"4bd4ff4d",
   854 => x"dbc21e75",
   855 => x"d7e849ec",
   856 => x"7086c487",
   857 => x"ccc40298",
   858 => x"48a6c487",
   859 => x"bff5ddc1",
   860 => x"fb497578",
   861 => x"d0ff87ef",
   862 => x"c178c548",
   863 => x"4ac07bd6",
   864 => x"1149a275",
   865 => x"cb82c17b",
   866 => x"f304aab7",
   867 => x"c34acc87",
   868 => x"82c17bff",
   869 => x"aab7e0c0",
   870 => x"ff87f404",
   871 => x"78c448d0",
   872 => x"c57bffc3",
   873 => x"7bd3c178",
   874 => x"78c47bc1",
   875 => x"b7c04866",
   876 => x"f0c206a8",
   877 => x"f4dbc287",
   878 => x"66c44cbf",
   879 => x"c8887448",
   880 => x"9c7458a6",
   881 => x"87f9c102",
   882 => x"7ef6cec2",
   883 => x"8c4dc0c8",
   884 => x"03acb7c0",
   885 => x"c0c887c6",
   886 => x"4cc04da4",
   887 => x"97e7dbc2",
   888 => x"99d049bf",
   889 => x"c087d102",
   890 => x"ecdbc21e",
   891 => x"87fbea49",
   892 => x"497086c4",
   893 => x"87eec04a",
   894 => x"1ef6cec2",
   895 => x"49ecdbc2",
   896 => x"c487e8ea",
   897 => x"4a497086",
   898 => x"c848d0ff",
   899 => x"d4c178c5",
   900 => x"bf976e7b",
   901 => x"c1486e7b",
   902 => x"c17e7080",
   903 => x"f0ff058d",
   904 => x"48d0ff87",
   905 => x"9a7278c4",
   906 => x"c087c505",
   907 => x"87c7c148",
   908 => x"dbc21ec1",
   909 => x"d8e849ec",
   910 => x"7486c487",
   911 => x"c7fe059c",
   912 => x"4866c487",
   913 => x"06a8b7c0",
   914 => x"dbc287d1",
   915 => x"78c048ec",
   916 => x"78c080d0",
   917 => x"dbc280f4",
   918 => x"c478bff8",
   919 => x"b7c04866",
   920 => x"d0fd01a8",
   921 => x"48d0ff87",
   922 => x"d3c178c5",
   923 => x"c47bc07b",
   924 => x"c248c178",
   925 => x"f848c087",
   926 => x"264d268e",
   927 => x"264b264c",
   928 => x"5b5e0e4f",
   929 => x"1e0e5d5c",
   930 => x"4cc04b71",
   931 => x"c004ab4d",
   932 => x"f2c087e8",
   933 => x"9d751edd",
   934 => x"c087c402",
   935 => x"c187c24a",
   936 => x"eb49724a",
   937 => x"86c487ea",
   938 => x"84c17e70",
   939 => x"87c2056e",
   940 => x"85c14c73",
   941 => x"ff06ac73",
   942 => x"486e87d8",
   943 => x"87f9fe26",
   944 => x"c44a711e",
   945 => x"87c50566",
   946 => x"fef94972",
   947 => x"0e4f2687",
   948 => x"5d5c5b5e",
   949 => x"4c711e0e",
   950 => x"c291de49",
   951 => x"714dd4dc",
   952 => x"026d9785",
   953 => x"c287dcc1",
   954 => x"4abfc0dc",
   955 => x"49728274",
   956 => x"7087cefe",
   957 => x"c0026e7e",
   958 => x"dcc287f2",
   959 => x"4a6e4bc8",
   960 => x"c6ff49cb",
   961 => x"4b7487e2",
   962 => x"dec193cb",
   963 => x"83c483c7",
   964 => x"7bc7fdc0",
   965 => x"c1c14974",
   966 => x"7b7587e7",
   967 => x"97f4ddc1",
   968 => x"c21e49bf",
   969 => x"fe49c8dc",
   970 => x"86c487d6",
   971 => x"c1c14974",
   972 => x"49c087cf",
   973 => x"87eec2c1",
   974 => x"48e8dbc2",
   975 => x"49c178c0",
   976 => x"2687d9dd",
   977 => x"4c87f2fc",
   978 => x"6964616f",
   979 => x"2e2e676e",
   980 => x"5e0e002e",
   981 => x"710e5c5b",
   982 => x"dcc24a4b",
   983 => x"7282bfc0",
   984 => x"87ddfc49",
   985 => x"029c4c70",
   986 => x"e74987c4",
   987 => x"dcc287ea",
   988 => x"78c048c0",
   989 => x"e3dc49c1",
   990 => x"87fffb87",
   991 => x"5c5b5e0e",
   992 => x"86f40e5d",
   993 => x"4df6cec2",
   994 => x"a6c44cc0",
   995 => x"c278c048",
   996 => x"49bfc0dc",
   997 => x"c106a9c0",
   998 => x"cec287c1",
   999 => x"029848f6",
  1000 => x"c087f8c0",
  1001 => x"c81eddf2",
  1002 => x"87c70266",
  1003 => x"c048a6c4",
  1004 => x"c487c578",
  1005 => x"78c148a6",
  1006 => x"e74966c4",
  1007 => x"86c487d2",
  1008 => x"84c14d70",
  1009 => x"c14866c4",
  1010 => x"58a6c880",
  1011 => x"bfc0dcc2",
  1012 => x"c603ac49",
  1013 => x"059d7587",
  1014 => x"c087c8ff",
  1015 => x"029d754c",
  1016 => x"c087e0c3",
  1017 => x"c81eddf2",
  1018 => x"87c70266",
  1019 => x"c048a6cc",
  1020 => x"cc87c578",
  1021 => x"78c148a6",
  1022 => x"e64966cc",
  1023 => x"86c487d2",
  1024 => x"026e7e70",
  1025 => x"6e87e9c2",
  1026 => x"9781cb49",
  1027 => x"99d04969",
  1028 => x"87d6c102",
  1029 => x"4ad2fdc0",
  1030 => x"91cb4974",
  1031 => x"81c7dec1",
  1032 => x"81c87972",
  1033 => x"7451ffc3",
  1034 => x"c291de49",
  1035 => x"714dd4dc",
  1036 => x"97c1c285",
  1037 => x"49a5c17d",
  1038 => x"c251e0c0",
  1039 => x"bf97c6d7",
  1040 => x"c187d202",
  1041 => x"4ba5c284",
  1042 => x"4ac6d7c2",
  1043 => x"c1ff49db",
  1044 => x"dbc187d6",
  1045 => x"49a5cd87",
  1046 => x"84c151c0",
  1047 => x"6e4ba5c2",
  1048 => x"ff49cb4a",
  1049 => x"c187c1c1",
  1050 => x"fbc087c6",
  1051 => x"49744acf",
  1052 => x"dec191cb",
  1053 => x"797281c7",
  1054 => x"97c6d7c2",
  1055 => x"87d802bf",
  1056 => x"91de4974",
  1057 => x"dcc284c1",
  1058 => x"83714bd4",
  1059 => x"4ac6d7c2",
  1060 => x"c0ff49dd",
  1061 => x"87d887d2",
  1062 => x"93de4b74",
  1063 => x"83d4dcc2",
  1064 => x"c049a3cb",
  1065 => x"7384c151",
  1066 => x"49cb4a6e",
  1067 => x"87f8fffe",
  1068 => x"c14866c4",
  1069 => x"58a6c880",
  1070 => x"c003acc7",
  1071 => x"056e87c5",
  1072 => x"7487e0fc",
  1073 => x"f68ef448",
  1074 => x"731e87ef",
  1075 => x"494b711e",
  1076 => x"dec191cb",
  1077 => x"a1c881c7",
  1078 => x"f3ddc14a",
  1079 => x"c9501248",
  1080 => x"f5c04aa1",
  1081 => x"501248ca",
  1082 => x"ddc181ca",
  1083 => x"501148f4",
  1084 => x"97f4ddc1",
  1085 => x"c01e49bf",
  1086 => x"87c4f749",
  1087 => x"48e8dbc2",
  1088 => x"49c178de",
  1089 => x"2687d5d6",
  1090 => x"1e87f2f5",
  1091 => x"cb494a71",
  1092 => x"c7dec191",
  1093 => x"1181c881",
  1094 => x"ecdbc248",
  1095 => x"c0dcc258",
  1096 => x"c178c048",
  1097 => x"87f4d549",
  1098 => x"c01e4f26",
  1099 => x"f5fac049",
  1100 => x"1e4f2687",
  1101 => x"d2029971",
  1102 => x"dcdfc187",
  1103 => x"f750c048",
  1104 => x"cbc4c180",
  1105 => x"c0dec140",
  1106 => x"c187ce78",
  1107 => x"c148d8df",
  1108 => x"fc78f9dd",
  1109 => x"eac4c180",
  1110 => x"0e4f2678",
  1111 => x"0e5c5b5e",
  1112 => x"cb4a4c71",
  1113 => x"c7dec192",
  1114 => x"49a2c882",
  1115 => x"974ba2c9",
  1116 => x"971e4b6b",
  1117 => x"ca1e4969",
  1118 => x"c0491282",
  1119 => x"c087f0e5",
  1120 => x"87d8d449",
  1121 => x"f7c04974",
  1122 => x"8ef887f7",
  1123 => x"1e87ecf3",
  1124 => x"4b711e73",
  1125 => x"87c3ff49",
  1126 => x"fefe4973",
  1127 => x"87ddf387",
  1128 => x"711e731e",
  1129 => x"4aa3c64b",
  1130 => x"c187db02",
  1131 => x"87d6028a",
  1132 => x"dac1028a",
  1133 => x"c0028a87",
  1134 => x"028a87fc",
  1135 => x"8a87e1c0",
  1136 => x"c187cb02",
  1137 => x"49c787db",
  1138 => x"c187c0fd",
  1139 => x"dcc287de",
  1140 => x"c102bfc0",
  1141 => x"c14887cb",
  1142 => x"c4dcc288",
  1143 => x"87c1c158",
  1144 => x"bfc4dcc2",
  1145 => x"87f9c002",
  1146 => x"bfc0dcc2",
  1147 => x"c280c148",
  1148 => x"c058c4dc",
  1149 => x"dcc287eb",
  1150 => x"c649bfc0",
  1151 => x"c4dcc289",
  1152 => x"a9b7c059",
  1153 => x"c287da03",
  1154 => x"c048c0dc",
  1155 => x"c287d278",
  1156 => x"02bfc4dc",
  1157 => x"dcc287cb",
  1158 => x"c648bfc0",
  1159 => x"c4dcc280",
  1160 => x"d149c058",
  1161 => x"497387f6",
  1162 => x"87d5f5c0",
  1163 => x"0e87cef1",
  1164 => x"5d5c5b5e",
  1165 => x"86d0ff0e",
  1166 => x"c859a6dc",
  1167 => x"78c048a6",
  1168 => x"c4c180c4",
  1169 => x"80c47866",
  1170 => x"80c478c1",
  1171 => x"dcc278c1",
  1172 => x"78c148c4",
  1173 => x"bfe8dbc2",
  1174 => x"05a8de48",
  1175 => x"dbf487cb",
  1176 => x"cc497087",
  1177 => x"f2cf59a6",
  1178 => x"87e8e487",
  1179 => x"e487cae5",
  1180 => x"4c7087d7",
  1181 => x"02acfbc0",
  1182 => x"d887fbc1",
  1183 => x"edc10566",
  1184 => x"66c0c187",
  1185 => x"6a82c44a",
  1186 => x"c11e727e",
  1187 => x"c448d0da",
  1188 => x"a1c84966",
  1189 => x"7141204a",
  1190 => x"87f905aa",
  1191 => x"4a265110",
  1192 => x"4866c0c1",
  1193 => x"78cac3c1",
  1194 => x"81c7496a",
  1195 => x"c0c15174",
  1196 => x"81c84966",
  1197 => x"c0c151c1",
  1198 => x"81c94966",
  1199 => x"c0c151c0",
  1200 => x"81ca4966",
  1201 => x"1ec151c0",
  1202 => x"496a1ed8",
  1203 => x"fce381c8",
  1204 => x"c186c887",
  1205 => x"c04866c4",
  1206 => x"87c701a8",
  1207 => x"c148a6c8",
  1208 => x"c187ce78",
  1209 => x"c14866c4",
  1210 => x"58a6d088",
  1211 => x"c8e387c3",
  1212 => x"48a6d087",
  1213 => x"9c7478c2",
  1214 => x"87dbcd02",
  1215 => x"c14866c8",
  1216 => x"03a866c8",
  1217 => x"dc87d0cd",
  1218 => x"78c048a6",
  1219 => x"78c080e8",
  1220 => x"7087f6e1",
  1221 => x"acd0c14c",
  1222 => x"87d7c205",
  1223 => x"e47e66c4",
  1224 => x"497087da",
  1225 => x"e159a6c8",
  1226 => x"4c7087df",
  1227 => x"05acecc0",
  1228 => x"c887ebc1",
  1229 => x"91cb4966",
  1230 => x"8166c0c1",
  1231 => x"6a4aa1c4",
  1232 => x"4aa1c84d",
  1233 => x"c15266c4",
  1234 => x"e079cbc4",
  1235 => x"4c7087fb",
  1236 => x"87d8029c",
  1237 => x"02acfbc0",
  1238 => x"557487d2",
  1239 => x"7087eae0",
  1240 => x"c7029c4c",
  1241 => x"acfbc087",
  1242 => x"87eeff05",
  1243 => x"c255e0c0",
  1244 => x"97c055c1",
  1245 => x"4966d87d",
  1246 => x"db05a96e",
  1247 => x"4866c887",
  1248 => x"04a866cc",
  1249 => x"66c887ca",
  1250 => x"cc80c148",
  1251 => x"87c858a6",
  1252 => x"c14866cc",
  1253 => x"58a6d088",
  1254 => x"87eddfff",
  1255 => x"d0c14c70",
  1256 => x"87c805ac",
  1257 => x"c14866d4",
  1258 => x"58a6d880",
  1259 => x"02acd0c1",
  1260 => x"c087e9fd",
  1261 => x"d848a6e0",
  1262 => x"66c47866",
  1263 => x"66e0c048",
  1264 => x"e4c905a8",
  1265 => x"a6e4c087",
  1266 => x"c478c048",
  1267 => x"7478c080",
  1268 => x"88fbc048",
  1269 => x"026e7e70",
  1270 => x"6e87e7c8",
  1271 => x"7088cb48",
  1272 => x"c1026e7e",
  1273 => x"486e87cd",
  1274 => x"7e7088c9",
  1275 => x"e9c3026e",
  1276 => x"c4486e87",
  1277 => x"6e7e7088",
  1278 => x"6e87ce02",
  1279 => x"7088c148",
  1280 => x"c3026e7e",
  1281 => x"f3c787d4",
  1282 => x"48a6dc87",
  1283 => x"ff78f0c0",
  1284 => x"7087f6dd",
  1285 => x"acecc04c",
  1286 => x"87c4c002",
  1287 => x"5ca6e0c0",
  1288 => x"02acecc0",
  1289 => x"ddff87cd",
  1290 => x"4c7087df",
  1291 => x"05acecc0",
  1292 => x"c087f3ff",
  1293 => x"c002acec",
  1294 => x"ddff87c4",
  1295 => x"1ec087cb",
  1296 => x"66d01eca",
  1297 => x"c191cb49",
  1298 => x"714866c8",
  1299 => x"58a6cc80",
  1300 => x"c44866c8",
  1301 => x"58a6d080",
  1302 => x"49bf66cc",
  1303 => x"87edddff",
  1304 => x"1ede1ec1",
  1305 => x"49bf66d4",
  1306 => x"87e1ddff",
  1307 => x"497086d0",
  1308 => x"c08909c0",
  1309 => x"c059a6ec",
  1310 => x"c04866e8",
  1311 => x"eec006a8",
  1312 => x"66e8c087",
  1313 => x"03a8dd48",
  1314 => x"c487e4c0",
  1315 => x"c049bf66",
  1316 => x"c08166e8",
  1317 => x"e8c051e0",
  1318 => x"81c14966",
  1319 => x"81bf66c4",
  1320 => x"c051c1c2",
  1321 => x"c24966e8",
  1322 => x"bf66c481",
  1323 => x"6e51c081",
  1324 => x"cac3c148",
  1325 => x"c8496e78",
  1326 => x"5166d081",
  1327 => x"81c9496e",
  1328 => x"6e5166d4",
  1329 => x"dc81ca49",
  1330 => x"66d05166",
  1331 => x"d480c148",
  1332 => x"d84858a6",
  1333 => x"c478c180",
  1334 => x"ddff87e8",
  1335 => x"497087de",
  1336 => x"59a6ecc0",
  1337 => x"87d4ddff",
  1338 => x"e0c04970",
  1339 => x"66dc59a6",
  1340 => x"a8ecc048",
  1341 => x"87cac005",
  1342 => x"c048a6dc",
  1343 => x"c07866e8",
  1344 => x"daff87c4",
  1345 => x"66c887c3",
  1346 => x"c191cb49",
  1347 => x"714866c0",
  1348 => x"6e7e7080",
  1349 => x"6e82c84a",
  1350 => x"c081ca49",
  1351 => x"dc5166e8",
  1352 => x"81c14966",
  1353 => x"8966e8c0",
  1354 => x"307148c1",
  1355 => x"89c14970",
  1356 => x"c27a9771",
  1357 => x"49bff0df",
  1358 => x"2966e8c0",
  1359 => x"484a6a97",
  1360 => x"f0c09871",
  1361 => x"496e58a6",
  1362 => x"4d6981c4",
  1363 => x"4866e0c0",
  1364 => x"02a866c4",
  1365 => x"c487c8c0",
  1366 => x"78c048a6",
  1367 => x"c487c5c0",
  1368 => x"78c148a6",
  1369 => x"c01e66c4",
  1370 => x"49751ee0",
  1371 => x"87ddd9ff",
  1372 => x"4c7086c8",
  1373 => x"06acb7c0",
  1374 => x"7487d4c1",
  1375 => x"49e0c085",
  1376 => x"4b758974",
  1377 => x"4ad9dac1",
  1378 => x"dbecfe71",
  1379 => x"c085c287",
  1380 => x"c14866e4",
  1381 => x"a6e8c080",
  1382 => x"66ecc058",
  1383 => x"7081c149",
  1384 => x"c8c002a9",
  1385 => x"48a6c487",
  1386 => x"c5c078c0",
  1387 => x"48a6c487",
  1388 => x"66c478c1",
  1389 => x"49a4c21e",
  1390 => x"7148e0c0",
  1391 => x"1e497088",
  1392 => x"d8ff4975",
  1393 => x"86c887c7",
  1394 => x"01a8b7c0",
  1395 => x"c087c0ff",
  1396 => x"c00266e4",
  1397 => x"496e87d1",
  1398 => x"e4c081c9",
  1399 => x"486e5166",
  1400 => x"78dbc5c1",
  1401 => x"6e87ccc0",
  1402 => x"c281c949",
  1403 => x"c1486e51",
  1404 => x"c078cfc6",
  1405 => x"c148a6e8",
  1406 => x"87c6c078",
  1407 => x"87f9d6ff",
  1408 => x"e8c04c70",
  1409 => x"f5c00266",
  1410 => x"4866c887",
  1411 => x"04a866cc",
  1412 => x"c887cbc0",
  1413 => x"80c14866",
  1414 => x"c058a6cc",
  1415 => x"66cc87e0",
  1416 => x"d088c148",
  1417 => x"d5c058a6",
  1418 => x"acc6c187",
  1419 => x"87c8c005",
  1420 => x"c14866d0",
  1421 => x"58a6d480",
  1422 => x"87fdd5ff",
  1423 => x"66d44c70",
  1424 => x"d880c148",
  1425 => x"9c7458a6",
  1426 => x"87cbc002",
  1427 => x"c14866c8",
  1428 => x"04a866c8",
  1429 => x"ff87f0f2",
  1430 => x"c887d5d5",
  1431 => x"a8c74866",
  1432 => x"87e5c003",
  1433 => x"48c4dcc2",
  1434 => x"66c878c0",
  1435 => x"c191cb49",
  1436 => x"c48166c0",
  1437 => x"4a6a4aa1",
  1438 => x"c87952c0",
  1439 => x"80c14866",
  1440 => x"c758a6cc",
  1441 => x"dbff04a8",
  1442 => x"8ed0ff87",
  1443 => x"87e9dfff",
  1444 => x"64616f4c",
  1445 => x"202e2a20",
  1446 => x"00203a00",
  1447 => x"711e731e",
  1448 => x"c6029b4b",
  1449 => x"c0dcc287",
  1450 => x"c778c048",
  1451 => x"c0dcc21e",
  1452 => x"c11e49bf",
  1453 => x"c21ec7de",
  1454 => x"49bfe8db",
  1455 => x"cc87f0ed",
  1456 => x"e8dbc286",
  1457 => x"eae949bf",
  1458 => x"029b7387",
  1459 => x"dec187c8",
  1460 => x"e3c049c7",
  1461 => x"deff87fd",
  1462 => x"c11e87e3",
  1463 => x"c048f3dd",
  1464 => x"eadfc150",
  1465 => x"d9ff49bf",
  1466 => x"48c087e1",
  1467 => x"c71e4f26",
  1468 => x"49c187df",
  1469 => x"fe87e5fe",
  1470 => x"7087eeee",
  1471 => x"87cd0298",
  1472 => x"87c7f6fe",
  1473 => x"c4029870",
  1474 => x"c24ac187",
  1475 => x"724ac087",
  1476 => x"87ce059a",
  1477 => x"dcc11ec0",
  1478 => x"efc049fe",
  1479 => x"86c487c3",
  1480 => x"1ec087fe",
  1481 => x"49c9ddc1",
  1482 => x"87f5eec0",
  1483 => x"e9fe1ec0",
  1484 => x"c0497087",
  1485 => x"c387eaee",
  1486 => x"8ef887d6",
  1487 => x"44534f26",
  1488 => x"69616620",
  1489 => x"2e64656c",
  1490 => x"6f6f4200",
  1491 => x"676e6974",
  1492 => x"002e2e2e",
  1493 => x"d6e6c01e",
  1494 => x"2687fa87",
  1495 => x"dcc21e4f",
  1496 => x"78c048c0",
  1497 => x"48e8dbc2",
  1498 => x"c1fe78c0",
  1499 => x"c087e587",
  1500 => x"004f2648",
  1501 => x"00000100",
  1502 => x"45208000",
  1503 => x"00746978",
  1504 => x"61422080",
  1505 => x"0b006b63",
  1506 => x"14000011",
  1507 => x"00000027",
  1508 => x"110b0000",
  1509 => x"27320000",
  1510 => x"00000000",
  1511 => x"00110b00",
  1512 => x"00275000",
  1513 => x"00000000",
  1514 => x"0000110b",
  1515 => x"0000276e",
  1516 => x"0b000000",
  1517 => x"8c000011",
  1518 => x"00000027",
  1519 => x"110b0000",
  1520 => x"27aa0000",
  1521 => x"00000000",
  1522 => x"00110b00",
  1523 => x"0027c800",
  1524 => x"00000000",
  1525 => x"0000110b",
  1526 => x"00000000",
  1527 => x"a0000000",
  1528 => x"00000011",
  1529 => x"00000000",
  1530 => x"17ee0000",
  1531 => x"4f420000",
  1532 => x"2020544f",
  1533 => x"4f522020",
  1534 => x"fe1e004d",
  1535 => x"78c048f0",
  1536 => x"097909cd",
  1537 => x"1e1e4f26",
  1538 => x"7ebff0fe",
  1539 => x"4f262648",
  1540 => x"48f0fe1e",
  1541 => x"4f2678c1",
  1542 => x"48f0fe1e",
  1543 => x"4f2678c0",
  1544 => x"c04a711e",
  1545 => x"4f265252",
  1546 => x"5c5b5e0e",
  1547 => x"86f40e5d",
  1548 => x"6d974d71",
  1549 => x"4ca5c17e",
  1550 => x"c8486c97",
  1551 => x"486e58a6",
  1552 => x"05a866c4",
  1553 => x"48ff87c5",
  1554 => x"ff87e6c0",
  1555 => x"a5c287ca",
  1556 => x"4b6c9749",
  1557 => x"974ba371",
  1558 => x"6c974b6b",
  1559 => x"c1486e7e",
  1560 => x"58a6c880",
  1561 => x"a6cc98c7",
  1562 => x"7c977058",
  1563 => x"7387e1fe",
  1564 => x"268ef448",
  1565 => x"264c264d",
  1566 => x"0e4f264b",
  1567 => x"0e5c5b5e",
  1568 => x"4c7186f4",
  1569 => x"c34a66d8",
  1570 => x"a4c29aff",
  1571 => x"496c974b",
  1572 => x"7249a173",
  1573 => x"7e6c9751",
  1574 => x"80c1486e",
  1575 => x"c758a6c8",
  1576 => x"58a6cc98",
  1577 => x"8ef45470",
  1578 => x"1e87caff",
  1579 => x"87e8fd1e",
  1580 => x"494abfe0",
  1581 => x"99c0e0c0",
  1582 => x"7287cb02",
  1583 => x"e6dfc21e",
  1584 => x"87f7fe49",
  1585 => x"fdfc86c4",
  1586 => x"fd7e7087",
  1587 => x"262687c2",
  1588 => x"dfc21e4f",
  1589 => x"c7fd49e6",
  1590 => x"ebe2c187",
  1591 => x"87dafc49",
  1592 => x"2687c7c4",
  1593 => x"d0ff1e4f",
  1594 => x"78e1c848",
  1595 => x"c548d4ff",
  1596 => x"0266c478",
  1597 => x"e0c387c3",
  1598 => x"0266c878",
  1599 => x"d4ff87c6",
  1600 => x"78f0c348",
  1601 => x"7148d4ff",
  1602 => x"48d0ff78",
  1603 => x"c078e1c8",
  1604 => x"4f2678e0",
  1605 => x"5c5b5e0e",
  1606 => x"c24c710e",
  1607 => x"fc49e6df",
  1608 => x"4a7087c6",
  1609 => x"04aab7c0",
  1610 => x"c387e2c2",
  1611 => x"c905aaf0",
  1612 => x"d9e7c187",
  1613 => x"c278c148",
  1614 => x"e0c387c3",
  1615 => x"87c905aa",
  1616 => x"48dde7c1",
  1617 => x"f4c178c1",
  1618 => x"dde7c187",
  1619 => x"87c602bf",
  1620 => x"4ba2c0c2",
  1621 => x"4b7287c2",
  1622 => x"d1059c74",
  1623 => x"d9e7c187",
  1624 => x"e7c11ebf",
  1625 => x"721ebfdd",
  1626 => x"87f9fd49",
  1627 => x"e7c186c8",
  1628 => x"c002bfd9",
  1629 => x"497387e0",
  1630 => x"9129b7c4",
  1631 => x"81f9e8c1",
  1632 => x"9acf4a73",
  1633 => x"48c192c2",
  1634 => x"4a703072",
  1635 => x"4872baff",
  1636 => x"79709869",
  1637 => x"497387db",
  1638 => x"9129b7c4",
  1639 => x"81f9e8c1",
  1640 => x"9acf4a73",
  1641 => x"48c392c2",
  1642 => x"4a703072",
  1643 => x"70b06948",
  1644 => x"dde7c179",
  1645 => x"c178c048",
  1646 => x"c048d9e7",
  1647 => x"e6dfc278",
  1648 => x"87e4f949",
  1649 => x"b7c04a70",
  1650 => x"defd03aa",
  1651 => x"c248c087",
  1652 => x"264d2687",
  1653 => x"264b264c",
  1654 => x"0000004f",
  1655 => x"00000000",
  1656 => x"4a711e00",
  1657 => x"87ecfc49",
  1658 => x"c01e4f26",
  1659 => x"c449724a",
  1660 => x"f9e8c191",
  1661 => x"c179c081",
  1662 => x"aab7d082",
  1663 => x"2687ee04",
  1664 => x"5b5e0e4f",
  1665 => x"710e5d5c",
  1666 => x"87ccf84d",
  1667 => x"b7c44a75",
  1668 => x"e8c1922a",
  1669 => x"4c7582f9",
  1670 => x"94c29ccf",
  1671 => x"744b496a",
  1672 => x"c29bc32b",
  1673 => x"70307448",
  1674 => x"74bcff4c",
  1675 => x"70987148",
  1676 => x"87dcf77a",
  1677 => x"d8fe4873",
  1678 => x"00000087",
  1679 => x"00000000",
  1680 => x"00000000",
  1681 => x"00000000",
  1682 => x"00000000",
  1683 => x"00000000",
  1684 => x"00000000",
  1685 => x"00000000",
  1686 => x"00000000",
  1687 => x"00000000",
  1688 => x"00000000",
  1689 => x"00000000",
  1690 => x"00000000",
  1691 => x"00000000",
  1692 => x"00000000",
  1693 => x"00000000",
  1694 => x"d0ff1e00",
  1695 => x"78e1c848",
  1696 => x"d4ff4871",
  1697 => x"66c47808",
  1698 => x"08d4ff48",
  1699 => x"1e4f2678",
  1700 => x"66c44a71",
  1701 => x"49721e49",
  1702 => x"ff87deff",
  1703 => x"e0c048d0",
  1704 => x"4f262678",
  1705 => x"711e731e",
  1706 => x"4966c84b",
  1707 => x"c14a731e",
  1708 => x"ff49a2e0",
  1709 => x"c42687d9",
  1710 => x"264d2687",
  1711 => x"264b264c",
  1712 => x"d4ff1e4f",
  1713 => x"7affc34a",
  1714 => x"c048d0ff",
  1715 => x"7ade78e1",
  1716 => x"bff0dfc2",
  1717 => x"c848497a",
  1718 => x"717a7028",
  1719 => x"7028d048",
  1720 => x"d848717a",
  1721 => x"ff7a7028",
  1722 => x"e0c048d0",
  1723 => x"0e4f2678",
  1724 => x"5d5c5b5e",
  1725 => x"c24c710e",
  1726 => x"4dbff0df",
  1727 => x"d02b744b",
  1728 => x"83c19b66",
  1729 => x"04ab66d4",
  1730 => x"4bc087c2",
  1731 => x"66d04a74",
  1732 => x"ff317249",
  1733 => x"739975b9",
  1734 => x"70307248",
  1735 => x"b071484a",
  1736 => x"58f4dfc2",
  1737 => x"2687dafe",
  1738 => x"264c264d",
  1739 => x"1e4f264b",
  1740 => x"c848d0ff",
  1741 => x"487178c9",
  1742 => x"7808d4ff",
  1743 => x"711e4f26",
  1744 => x"87eb494a",
  1745 => x"c848d0ff",
  1746 => x"1e4f2678",
  1747 => x"4b711e73",
  1748 => x"bfc0e0c2",
  1749 => x"c287c302",
  1750 => x"d0ff87eb",
  1751 => x"78c9c848",
  1752 => x"e0c04973",
  1753 => x"48d4ffb1",
  1754 => x"dfc27871",
  1755 => x"78c048f4",
  1756 => x"c50266c8",
  1757 => x"49ffc387",
  1758 => x"49c087c2",
  1759 => x"59fcdfc2",
  1760 => x"c60266cc",
  1761 => x"d5d5c587",
  1762 => x"cf87c44a",
  1763 => x"c24affff",
  1764 => x"c25ac0e0",
  1765 => x"c148c0e0",
  1766 => x"2687c478",
  1767 => x"264c264d",
  1768 => x"0e4f264b",
  1769 => x"5d5c5b5e",
  1770 => x"c24a710e",
  1771 => x"4cbffcdf",
  1772 => x"cb029a72",
  1773 => x"91c84987",
  1774 => x"4bc1edc1",
  1775 => x"87c48371",
  1776 => x"4bc1f1c1",
  1777 => x"49134dc0",
  1778 => x"dfc29974",
  1779 => x"ffb9bff8",
  1780 => x"787148d4",
  1781 => x"852cb7c1",
  1782 => x"04adb7c8",
  1783 => x"dfc287e8",
  1784 => x"c848bff4",
  1785 => x"f8dfc280",
  1786 => x"87effe58",
  1787 => x"711e731e",
  1788 => x"9a4a134b",
  1789 => x"7287cb02",
  1790 => x"87e7fe49",
  1791 => x"059a4a13",
  1792 => x"dafe87f5",
  1793 => x"dfc21e87",
  1794 => x"c249bff4",
  1795 => x"c148f4df",
  1796 => x"c0c478a1",
  1797 => x"db03a9b7",
  1798 => x"48d4ff87",
  1799 => x"bff8dfc2",
  1800 => x"f4dfc278",
  1801 => x"dfc249bf",
  1802 => x"a1c148f4",
  1803 => x"b7c0c478",
  1804 => x"87e504a9",
  1805 => x"c848d0ff",
  1806 => x"c0e0c278",
  1807 => x"2678c048",
  1808 => x"0000004f",
  1809 => x"00000000",
  1810 => x"00000000",
  1811 => x"00005f5f",
  1812 => x"03030000",
  1813 => x"00030300",
  1814 => x"7f7f1400",
  1815 => x"147f7f14",
  1816 => x"2e240000",
  1817 => x"123a6b6b",
  1818 => x"366a4c00",
  1819 => x"32566c18",
  1820 => x"4f7e3000",
  1821 => x"683a7759",
  1822 => x"04000040",
  1823 => x"00000307",
  1824 => x"1c000000",
  1825 => x"0041633e",
  1826 => x"41000000",
  1827 => x"001c3e63",
  1828 => x"3e2a0800",
  1829 => x"2a3e1c1c",
  1830 => x"08080008",
  1831 => x"08083e3e",
  1832 => x"80000000",
  1833 => x"000060e0",
  1834 => x"08080000",
  1835 => x"08080808",
  1836 => x"00000000",
  1837 => x"00006060",
  1838 => x"30604000",
  1839 => x"03060c18",
  1840 => x"7f3e0001",
  1841 => x"3e7f4d59",
  1842 => x"06040000",
  1843 => x"00007f7f",
  1844 => x"63420000",
  1845 => x"464f5971",
  1846 => x"63220000",
  1847 => x"367f4949",
  1848 => x"161c1800",
  1849 => x"107f7f13",
  1850 => x"67270000",
  1851 => x"397d4545",
  1852 => x"7e3c0000",
  1853 => x"3079494b",
  1854 => x"01010000",
  1855 => x"070f7971",
  1856 => x"7f360000",
  1857 => x"367f4949",
  1858 => x"4f060000",
  1859 => x"1e3f6949",
  1860 => x"00000000",
  1861 => x"00006666",
  1862 => x"80000000",
  1863 => x"000066e6",
  1864 => x"08080000",
  1865 => x"22221414",
  1866 => x"14140000",
  1867 => x"14141414",
  1868 => x"22220000",
  1869 => x"08081414",
  1870 => x"03020000",
  1871 => x"060f5951",
  1872 => x"417f3e00",
  1873 => x"1e1f555d",
  1874 => x"7f7e0000",
  1875 => x"7e7f0909",
  1876 => x"7f7f0000",
  1877 => x"367f4949",
  1878 => x"3e1c0000",
  1879 => x"41414163",
  1880 => x"7f7f0000",
  1881 => x"1c3e6341",
  1882 => x"7f7f0000",
  1883 => x"41414949",
  1884 => x"7f7f0000",
  1885 => x"01010909",
  1886 => x"7f3e0000",
  1887 => x"7a7b4941",
  1888 => x"7f7f0000",
  1889 => x"7f7f0808",
  1890 => x"41000000",
  1891 => x"00417f7f",
  1892 => x"60200000",
  1893 => x"3f7f4040",
  1894 => x"087f7f00",
  1895 => x"4163361c",
  1896 => x"7f7f0000",
  1897 => x"40404040",
  1898 => x"067f7f00",
  1899 => x"7f7f060c",
  1900 => x"067f7f00",
  1901 => x"7f7f180c",
  1902 => x"7f3e0000",
  1903 => x"3e7f4141",
  1904 => x"7f7f0000",
  1905 => x"060f0909",
  1906 => x"417f3e00",
  1907 => x"407e7f61",
  1908 => x"7f7f0000",
  1909 => x"667f1909",
  1910 => x"6f260000",
  1911 => x"327b594d",
  1912 => x"01010000",
  1913 => x"01017f7f",
  1914 => x"7f3f0000",
  1915 => x"3f7f4040",
  1916 => x"3f0f0000",
  1917 => x"0f3f7070",
  1918 => x"307f7f00",
  1919 => x"7f7f3018",
  1920 => x"36634100",
  1921 => x"63361c1c",
  1922 => x"06030141",
  1923 => x"03067c7c",
  1924 => x"59716101",
  1925 => x"4143474d",
  1926 => x"7f000000",
  1927 => x"0041417f",
  1928 => x"06030100",
  1929 => x"6030180c",
  1930 => x"41000040",
  1931 => x"007f7f41",
  1932 => x"060c0800",
  1933 => x"080c0603",
  1934 => x"80808000",
  1935 => x"80808080",
  1936 => x"00000000",
  1937 => x"00040703",
  1938 => x"74200000",
  1939 => x"787c5454",
  1940 => x"7f7f0000",
  1941 => x"387c4444",
  1942 => x"7c380000",
  1943 => x"00444444",
  1944 => x"7c380000",
  1945 => x"7f7f4444",
  1946 => x"7c380000",
  1947 => x"185c5454",
  1948 => x"7e040000",
  1949 => x"0005057f",
  1950 => x"bc180000",
  1951 => x"7cfca4a4",
  1952 => x"7f7f0000",
  1953 => x"787c0404",
  1954 => x"00000000",
  1955 => x"00407d3d",
  1956 => x"80800000",
  1957 => x"007dfd80",
  1958 => x"7f7f0000",
  1959 => x"446c3810",
  1960 => x"00000000",
  1961 => x"00407f3f",
  1962 => x"0c7c7c00",
  1963 => x"787c0c18",
  1964 => x"7c7c0000",
  1965 => x"787c0404",
  1966 => x"7c380000",
  1967 => x"387c4444",
  1968 => x"fcfc0000",
  1969 => x"183c2424",
  1970 => x"3c180000",
  1971 => x"fcfc2424",
  1972 => x"7c7c0000",
  1973 => x"080c0404",
  1974 => x"5c480000",
  1975 => x"20745454",
  1976 => x"3f040000",
  1977 => x"0044447f",
  1978 => x"7c3c0000",
  1979 => x"7c7c4040",
  1980 => x"3c1c0000",
  1981 => x"1c3c6060",
  1982 => x"607c3c00",
  1983 => x"3c7c6030",
  1984 => x"386c4400",
  1985 => x"446c3810",
  1986 => x"bc1c0000",
  1987 => x"1c3c60e0",
  1988 => x"64440000",
  1989 => x"444c5c74",
  1990 => x"08080000",
  1991 => x"4141773e",
  1992 => x"00000000",
  1993 => x"00007f7f",
  1994 => x"41410000",
  1995 => x"08083e77",
  1996 => x"01010200",
  1997 => x"01020203",
  1998 => x"7f7f7f00",
  1999 => x"7f7f7f7f",
  2000 => x"1c080800",
  2001 => x"7f3e3e1c",
  2002 => x"3e7f7f7f",
  2003 => x"081c1c3e",
  2004 => x"18100008",
  2005 => x"10187c7c",
  2006 => x"30100000",
  2007 => x"10307c7c",
  2008 => x"60301000",
  2009 => x"061e7860",
  2010 => x"3c664200",
  2011 => x"42663c18",
  2012 => x"6a387800",
  2013 => x"386cc6c2",
  2014 => x"00006000",
  2015 => x"60000060",
  2016 => x"5b5e0e00",
  2017 => x"1e0e5d5c",
  2018 => x"e0c24c71",
  2019 => x"c04dbfd1",
  2020 => x"741ec04b",
  2021 => x"87c702ab",
  2022 => x"c048a6c4",
  2023 => x"c487c578",
  2024 => x"78c148a6",
  2025 => x"731e66c4",
  2026 => x"87dfee49",
  2027 => x"e0c086c8",
  2028 => x"87efef49",
  2029 => x"6a4aa5c4",
  2030 => x"87f0f049",
  2031 => x"cb87c6f1",
  2032 => x"c883c185",
  2033 => x"ff04abb7",
  2034 => x"262687c7",
  2035 => x"264c264d",
  2036 => x"1e4f264b",
  2037 => x"e0c24a71",
  2038 => x"e0c25ad5",
  2039 => x"78c748d5",
  2040 => x"87ddfe49",
  2041 => x"731e4f26",
  2042 => x"c04a711e",
  2043 => x"d303aab7",
  2044 => x"f6ccc287",
  2045 => x"87c405bf",
  2046 => x"87c24bc1",
  2047 => x"ccc24bc0",
  2048 => x"87c45bfa",
  2049 => x"5afaccc2",
  2050 => x"bff6ccc2",
  2051 => x"c19ac14a",
  2052 => x"ec49a2c0",
  2053 => x"48fc87e8",
  2054 => x"bff6ccc2",
  2055 => x"87effe78",
  2056 => x"c44a711e",
  2057 => x"49721e66",
  2058 => x"2687f9e9",
  2059 => x"c21e4f26",
  2060 => x"49bff6cc",
  2061 => x"c287eae6",
  2062 => x"e848c9e0",
  2063 => x"e0c278bf",
  2064 => x"bfec48c5",
  2065 => x"c9e0c278",
  2066 => x"c3494abf",
  2067 => x"b7c899ff",
  2068 => x"7148722a",
  2069 => x"d1e0c2b0",
  2070 => x"0e4f2658",
  2071 => x"5d5c5b5e",
  2072 => x"ff4b710e",
  2073 => x"e0c287c8",
  2074 => x"50c048c4",
  2075 => x"d0e64973",
  2076 => x"4c497087",
  2077 => x"eecb9cc2",
  2078 => x"87c2cb49",
  2079 => x"c24d4970",
  2080 => x"bf97c4e0",
  2081 => x"87e2c105",
  2082 => x"c24966d0",
  2083 => x"99bfcde0",
  2084 => x"d487d605",
  2085 => x"e0c24966",
  2086 => x"0599bfc5",
  2087 => x"497387cb",
  2088 => x"7087dee5",
  2089 => x"c1c10298",
  2090 => x"fe4cc187",
  2091 => x"497587c0",
  2092 => x"7087d7ca",
  2093 => x"87c60298",
  2094 => x"48c4e0c2",
  2095 => x"e0c250c1",
  2096 => x"05bf97c4",
  2097 => x"c287e3c0",
  2098 => x"49bfcde0",
  2099 => x"059966d0",
  2100 => x"c287d6ff",
  2101 => x"49bfc5e0",
  2102 => x"059966d4",
  2103 => x"7387caff",
  2104 => x"87dde449",
  2105 => x"fe059870",
  2106 => x"487487ff",
  2107 => x"0e87dcfb",
  2108 => x"5d5c5b5e",
  2109 => x"c086f40e",
  2110 => x"bfec4c4d",
  2111 => x"48a6c47e",
  2112 => x"bfd1e0c2",
  2113 => x"c01ec178",
  2114 => x"fd49c71e",
  2115 => x"86c887cd",
  2116 => x"cd029870",
  2117 => x"fb49ff87",
  2118 => x"dac187cc",
  2119 => x"87e1e349",
  2120 => x"e0c24dc1",
  2121 => x"02bf97c4",
  2122 => x"f6c887c3",
  2123 => x"c9e0c287",
  2124 => x"ccc24bbf",
  2125 => x"c005bff6",
  2126 => x"fdc387e9",
  2127 => x"87c1e349",
  2128 => x"e249fac3",
  2129 => x"497387fb",
  2130 => x"7199ffc3",
  2131 => x"fb49c01e",
  2132 => x"497387ce",
  2133 => x"7129b7c8",
  2134 => x"fb49c11e",
  2135 => x"86c887c2",
  2136 => x"c287f9c5",
  2137 => x"4bbfcde0",
  2138 => x"87dd029b",
  2139 => x"bff2ccc2",
  2140 => x"87d6c749",
  2141 => x"c4059870",
  2142 => x"d24bc087",
  2143 => x"49e0c287",
  2144 => x"c287fbc6",
  2145 => x"c658f6cc",
  2146 => x"f2ccc287",
  2147 => x"7378c048",
  2148 => x"0599c249",
  2149 => x"ebc387cd",
  2150 => x"87e5e149",
  2151 => x"99c24970",
  2152 => x"fb87c202",
  2153 => x"c149734c",
  2154 => x"87cd0599",
  2155 => x"e149f4c3",
  2156 => x"497087cf",
  2157 => x"c20299c2",
  2158 => x"734cfa87",
  2159 => x"0599c849",
  2160 => x"f5c387cd",
  2161 => x"87f9e049",
  2162 => x"99c24970",
  2163 => x"c287d402",
  2164 => x"02bfd5e0",
  2165 => x"c14887c9",
  2166 => x"d9e0c288",
  2167 => x"ff87c258",
  2168 => x"734dc14c",
  2169 => x"0599c449",
  2170 => x"f2c387cd",
  2171 => x"87d1e049",
  2172 => x"99c24970",
  2173 => x"c287db02",
  2174 => x"7ebfd5e0",
  2175 => x"a8b7c748",
  2176 => x"6e87cb03",
  2177 => x"c280c148",
  2178 => x"c058d9e0",
  2179 => x"4cfe87c2",
  2180 => x"fdc34dc1",
  2181 => x"e8dfff49",
  2182 => x"c2497087",
  2183 => x"87d50299",
  2184 => x"bfd5e0c2",
  2185 => x"87c9c002",
  2186 => x"48d5e0c2",
  2187 => x"c2c078c0",
  2188 => x"c14cfd87",
  2189 => x"49fac34d",
  2190 => x"87c5dfff",
  2191 => x"99c24970",
  2192 => x"c287d902",
  2193 => x"48bfd5e0",
  2194 => x"03a8b7c7",
  2195 => x"c287c9c0",
  2196 => x"c748d5e0",
  2197 => x"87c2c078",
  2198 => x"4dc14cfc",
  2199 => x"03acb7c0",
  2200 => x"c487d1c0",
  2201 => x"d8c14a66",
  2202 => x"c0026a82",
  2203 => x"4b6a87c6",
  2204 => x"0f734974",
  2205 => x"f0c31ec0",
  2206 => x"49dac11e",
  2207 => x"c887dcf7",
  2208 => x"02987086",
  2209 => x"c887e2c0",
  2210 => x"e0c248a6",
  2211 => x"c878bfd5",
  2212 => x"91cb4966",
  2213 => x"714866c4",
  2214 => x"6e7e7080",
  2215 => x"c8c002bf",
  2216 => x"4bbf6e87",
  2217 => x"734966c8",
  2218 => x"029d750f",
  2219 => x"c287c8c0",
  2220 => x"49bfd5e0",
  2221 => x"c287caf3",
  2222 => x"02bffacc",
  2223 => x"4987ddc0",
  2224 => x"7087c7c2",
  2225 => x"d3c00298",
  2226 => x"d5e0c287",
  2227 => x"f0f249bf",
  2228 => x"f449c087",
  2229 => x"ccc287d0",
  2230 => x"78c048fa",
  2231 => x"eaf38ef4",
  2232 => x"5b5e0e87",
  2233 => x"1e0e5d5c",
  2234 => x"e0c24c71",
  2235 => x"c149bfd1",
  2236 => x"c14da1cd",
  2237 => x"7e6981d1",
  2238 => x"cf029c74",
  2239 => x"4ba5c487",
  2240 => x"e0c27b74",
  2241 => x"f349bfd1",
  2242 => x"7b6e87c9",
  2243 => x"c4059c74",
  2244 => x"c24bc087",
  2245 => x"734bc187",
  2246 => x"87caf349",
  2247 => x"c70266d4",
  2248 => x"87da4987",
  2249 => x"87c24a70",
  2250 => x"ccc24ac0",
  2251 => x"f2265afe",
  2252 => x"000087d9",
  2253 => x"00000000",
  2254 => x"00000000",
  2255 => x"711e0000",
  2256 => x"bfc8ff4a",
  2257 => x"48a17249",
  2258 => x"ff1e4f26",
  2259 => x"fe89bfc8",
  2260 => x"c0c0c0c0",
  2261 => x"c401a9c0",
  2262 => x"c24ac087",
  2263 => x"724ac187",
  2264 => x"1e4f2648",
  2265 => x"bfcccec2",
  2266 => x"c2b9c149",
  2267 => x"ff59d0ce",
  2268 => x"ffc348d4",
  2269 => x"48d0ff78",
  2270 => x"ff78e1c0",
  2271 => x"78c148d4",
  2272 => x"787131c4",
  2273 => x"c048d0ff",
  2274 => x"4f2678e0",
  2275 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
