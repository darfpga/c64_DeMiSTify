library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0000417f",
     1 => x"40602000",
     2 => x"003f7f40",
     3 => x"1c087f7f",
     4 => x"00416336",
     5 => x"407f7f00",
     6 => x"00404040",
     7 => x"0c067f7f",
     8 => x"007f7f06",
     9 => x"0c067f7f",
    10 => x"007f7f18",
    11 => x"417f3e00",
    12 => x"003e7f41",
    13 => x"097f7f00",
    14 => x"00060f09",
    15 => x"61417f3e",
    16 => x"00407e7f",
    17 => x"097f7f00",
    18 => x"00667f19",
    19 => x"4d6f2600",
    20 => x"00327b59",
    21 => x"7f010100",
    22 => x"0001017f",
    23 => x"407f3f00",
    24 => x"003f7f40",
    25 => x"703f0f00",
    26 => x"000f3f70",
    27 => x"18307f7f",
    28 => x"007f7f30",
    29 => x"1c366341",
    30 => x"4163361c",
    31 => x"7c060301",
    32 => x"0103067c",
    33 => x"4d597161",
    34 => x"00414347",
    35 => x"7f7f0000",
    36 => x"00004141",
    37 => x"0c060301",
    38 => x"40603018",
    39 => x"41410000",
    40 => x"00007f7f",
    41 => x"03060c08",
    42 => x"00080c06",
    43 => x"80808080",
    44 => x"00808080",
    45 => x"03000000",
    46 => x"00000407",
    47 => x"54742000",
    48 => x"00787c54",
    49 => x"447f7f00",
    50 => x"00387c44",
    51 => x"447c3800",
    52 => x"00004444",
    53 => x"447c3800",
    54 => x"007f7f44",
    55 => x"547c3800",
    56 => x"00185c54",
    57 => x"7f7e0400",
    58 => x"00000505",
    59 => x"a4bc1800",
    60 => x"007cfca4",
    61 => x"047f7f00",
    62 => x"00787c04",
    63 => x"3d000000",
    64 => x"0000407d",
    65 => x"80808000",
    66 => x"00007dfd",
    67 => x"107f7f00",
    68 => x"00446c38",
    69 => x"3f000000",
    70 => x"0000407f",
    71 => x"180c7c7c",
    72 => x"00787c0c",
    73 => x"047c7c00",
    74 => x"00787c04",
    75 => x"447c3800",
    76 => x"00387c44",
    77 => x"24fcfc00",
    78 => x"00183c24",
    79 => x"243c1800",
    80 => x"00fcfc24",
    81 => x"047c7c00",
    82 => x"00080c04",
    83 => x"545c4800",
    84 => x"00207454",
    85 => x"7f3f0400",
    86 => x"00004444",
    87 => x"407c3c00",
    88 => x"007c7c40",
    89 => x"603c1c00",
    90 => x"001c3c60",
    91 => x"30607c3c",
    92 => x"003c7c60",
    93 => x"10386c44",
    94 => x"00446c38",
    95 => x"e0bc1c00",
    96 => x"001c3c60",
    97 => x"74644400",
    98 => x"00444c5c",
    99 => x"3e080800",
   100 => x"00414177",
   101 => x"7f000000",
   102 => x"0000007f",
   103 => x"77414100",
   104 => x"0008083e",
   105 => x"03010102",
   106 => x"00010202",
   107 => x"7f7f7f7f",
   108 => x"007f7f7f",
   109 => x"1c1c0808",
   110 => x"7f7f3e3e",
   111 => x"3e3e7f7f",
   112 => x"08081c1c",
   113 => x"7c181000",
   114 => x"0010187c",
   115 => x"7c301000",
   116 => x"0010307c",
   117 => x"60603010",
   118 => x"00061e78",
   119 => x"183c6642",
   120 => x"0042663c",
   121 => x"c26a3878",
   122 => x"00386cc6",
   123 => x"60000060",
   124 => x"00600000",
   125 => x"5c5b5e0e",
   126 => x"711e0e5d",
   127 => x"d9f1c24c",
   128 => x"4bc04dbf",
   129 => x"ab741ec0",
   130 => x"c487c702",
   131 => x"78c048a6",
   132 => x"a6c487c5",
   133 => x"c478c148",
   134 => x"49731e66",
   135 => x"c887dfee",
   136 => x"49e0c086",
   137 => x"c487efef",
   138 => x"496a4aa5",
   139 => x"f187f0f0",
   140 => x"85cb87c6",
   141 => x"b7c883c1",
   142 => x"c7ff04ab",
   143 => x"4d262687",
   144 => x"4b264c26",
   145 => x"711e4f26",
   146 => x"ddf1c24a",
   147 => x"ddf1c25a",
   148 => x"4978c748",
   149 => x"2687ddfe",
   150 => x"1e731e4f",
   151 => x"b7c04a71",
   152 => x"87d303aa",
   153 => x"bff3d6c2",
   154 => x"c187c405",
   155 => x"c087c24b",
   156 => x"f7d6c24b",
   157 => x"c287c45b",
   158 => x"c25af7d6",
   159 => x"4abff3d6",
   160 => x"c0c19ac1",
   161 => x"e8ec49a2",
   162 => x"c248fc87",
   163 => x"78bff3d6",
   164 => x"1e87effe",
   165 => x"66c44a71",
   166 => x"e649721e",
   167 => x"262687e2",
   168 => x"d6c21e4f",
   169 => x"e349bff3",
   170 => x"f1c287c4",
   171 => x"bfe848d1",
   172 => x"cdf1c278",
   173 => x"78bfec48",
   174 => x"bfd1f1c2",
   175 => x"ffc3494a",
   176 => x"2ab7c899",
   177 => x"b0714872",
   178 => x"58d9f1c2",
   179 => x"5e0e4f26",
   180 => x"0e5d5c5b",
   181 => x"c8ff4b71",
   182 => x"ccf1c287",
   183 => x"7350c048",
   184 => x"87eae249",
   185 => x"c24c4970",
   186 => x"49eecb9c",
   187 => x"7087cccb",
   188 => x"f1c24d49",
   189 => x"05bf97cc",
   190 => x"d087e2c1",
   191 => x"f1c24966",
   192 => x"0599bfd5",
   193 => x"66d487d6",
   194 => x"cdf1c249",
   195 => x"cb0599bf",
   196 => x"e1497387",
   197 => x"987087f8",
   198 => x"87c1c102",
   199 => x"c0fe4cc1",
   200 => x"ca497587",
   201 => x"987087e1",
   202 => x"c287c602",
   203 => x"c148ccf1",
   204 => x"ccf1c250",
   205 => x"c005bf97",
   206 => x"f1c287e3",
   207 => x"d049bfd5",
   208 => x"ff059966",
   209 => x"f1c287d6",
   210 => x"d449bfcd",
   211 => x"ff059966",
   212 => x"497387ca",
   213 => x"7087f7e0",
   214 => x"fffe0598",
   215 => x"fb487487",
   216 => x"5e0e87dc",
   217 => x"0e5d5c5b",
   218 => x"4dc086f4",
   219 => x"7ebfec4c",
   220 => x"c248a6c4",
   221 => x"78bfd9f1",
   222 => x"1ec01ec1",
   223 => x"cdfd49c7",
   224 => x"7086c887",
   225 => x"87ce0298",
   226 => x"ccfb49ff",
   227 => x"49dac187",
   228 => x"87fadfff",
   229 => x"f1c24dc1",
   230 => x"02bf97cc",
   231 => x"c4d087c3",
   232 => x"d1f1c287",
   233 => x"d6c24bbf",
   234 => x"c005bff3",
   235 => x"fdc387eb",
   236 => x"d9dfff49",
   237 => x"49fac387",
   238 => x"87d2dfff",
   239 => x"ffc34973",
   240 => x"c01e7199",
   241 => x"87cbfb49",
   242 => x"b7c84973",
   243 => x"c11e7129",
   244 => x"87fffa49",
   245 => x"c0c686c8",
   246 => x"d5f1c287",
   247 => x"029b4bbf",
   248 => x"d6c287dd",
   249 => x"c749bfef",
   250 => x"987087dd",
   251 => x"c087c405",
   252 => x"c287d24b",
   253 => x"c2c749e0",
   254 => x"f3d6c287",
   255 => x"c287c658",
   256 => x"c048efd6",
   257 => x"c2497378",
   258 => x"87ce0599",
   259 => x"ff49ebc3",
   260 => x"7087fbdd",
   261 => x"0299c249",
   262 => x"4cfb87c2",
   263 => x"99c14973",
   264 => x"c387ce05",
   265 => x"ddff49f4",
   266 => x"497087e4",
   267 => x"c20299c2",
   268 => x"734cfa87",
   269 => x"0599c849",
   270 => x"f5c387ce",
   271 => x"cdddff49",
   272 => x"c2497087",
   273 => x"87d50299",
   274 => x"bfddf1c2",
   275 => x"4887ca02",
   276 => x"f1c288c1",
   277 => x"c2c058e1",
   278 => x"c14cff87",
   279 => x"c449734d",
   280 => x"87ce0599",
   281 => x"ff49f2c3",
   282 => x"7087e3dc",
   283 => x"0299c249",
   284 => x"f1c287dc",
   285 => x"487ebfdd",
   286 => x"03a8b7c7",
   287 => x"6e87cbc0",
   288 => x"c280c148",
   289 => x"c058e1f1",
   290 => x"4cfe87c2",
   291 => x"fdc34dc1",
   292 => x"f9dbff49",
   293 => x"c2497087",
   294 => x"87d50299",
   295 => x"bfddf1c2",
   296 => x"87c9c002",
   297 => x"48ddf1c2",
   298 => x"c2c078c0",
   299 => x"c14cfd87",
   300 => x"49fac34d",
   301 => x"87d6dbff",
   302 => x"99c24970",
   303 => x"87d9c002",
   304 => x"bfddf1c2",
   305 => x"a8b7c748",
   306 => x"87c9c003",
   307 => x"48ddf1c2",
   308 => x"c2c078c7",
   309 => x"c14cfc87",
   310 => x"acb7c04d",
   311 => x"87d1c003",
   312 => x"c14a66c4",
   313 => x"026a82d8",
   314 => x"6a87c6c0",
   315 => x"7349744b",
   316 => x"c31ec00f",
   317 => x"dac11ef0",
   318 => x"87d2f749",
   319 => x"987086c8",
   320 => x"87e2c002",
   321 => x"c248a6c8",
   322 => x"78bfddf1",
   323 => x"cb4966c8",
   324 => x"4866c491",
   325 => x"7e708071",
   326 => x"c002bf6e",
   327 => x"bf6e87c8",
   328 => x"4966c84b",
   329 => x"9d750f73",
   330 => x"87c8c002",
   331 => x"bfddf1c2",
   332 => x"87c0f349",
   333 => x"bff7d6c2",
   334 => x"87ddc002",
   335 => x"87c7c249",
   336 => x"c0029870",
   337 => x"f1c287d3",
   338 => x"f249bfdd",
   339 => x"49c087e6",
   340 => x"c287c6f4",
   341 => x"c048f7d6",
   342 => x"f38ef478",
   343 => x"5e0e87e0",
   344 => x"0e5d5c5b",
   345 => x"c24c711e",
   346 => x"49bfd9f1",
   347 => x"4da1cdc1",
   348 => x"6981d1c1",
   349 => x"029c747e",
   350 => x"a5c487cf",
   351 => x"c27b744b",
   352 => x"49bfd9f1",
   353 => x"6e87fff2",
   354 => x"059c747b",
   355 => x"4bc087c4",
   356 => x"4bc187c2",
   357 => x"c0f34973",
   358 => x"0266d487",
   359 => x"da4987c7",
   360 => x"c24a7087",
   361 => x"c24ac087",
   362 => x"265afbd6",
   363 => x"0087cff2",
   364 => x"00000000",
   365 => x"00000000",
   366 => x"1e000000",
   367 => x"c8ff4a71",
   368 => x"a17249bf",
   369 => x"1e4f2648",
   370 => x"89bfc8ff",
   371 => x"c0c0c0fe",
   372 => x"01a9c0c0",
   373 => x"4ac087c4",
   374 => x"4ac187c2",
   375 => x"4f264872",
   376 => x"5c5b5e0e",
   377 => x"4b710e5d",
   378 => x"d04cd4ff",
   379 => x"78c04866",
   380 => x"d8ff49d6",
   381 => x"ffc387d0",
   382 => x"c3496c7c",
   383 => x"4d7199ff",
   384 => x"99f0c349",
   385 => x"05a9e0c1",
   386 => x"ffc387cb",
   387 => x"c3486c7c",
   388 => x"0866d098",
   389 => x"7cffc378",
   390 => x"c8494a6c",
   391 => x"7cffc331",
   392 => x"b2714a6c",
   393 => x"31c84972",
   394 => x"6c7cffc3",
   395 => x"72b2714a",
   396 => x"c331c849",
   397 => x"4a6c7cff",
   398 => x"d0ffb271",
   399 => x"78e0c048",
   400 => x"c2029b73",
   401 => x"757b7287",
   402 => x"264d2648",
   403 => x"264b264c",
   404 => x"4f261e4f",
   405 => x"5c5b5e0e",
   406 => x"7686f80e",
   407 => x"49a6c81e",
   408 => x"c487fdfd",
   409 => x"6e4b7086",
   410 => x"03a8c248",
   411 => x"7387f0c2",
   412 => x"9af0c34a",
   413 => x"02aad0c1",
   414 => x"e0c187c7",
   415 => x"dec205aa",
   416 => x"c8497387",
   417 => x"87c30299",
   418 => x"7387c6ff",
   419 => x"c29cc34c",
   420 => x"c2c105ac",
   421 => x"4966c487",
   422 => x"1e7131c9",
   423 => x"d44a66c4",
   424 => x"e1f1c292",
   425 => x"fe817249",
   426 => x"d887e7cc",
   427 => x"d5d5ff49",
   428 => x"1ec0c887",
   429 => x"49fadfc2",
   430 => x"87e3e8fd",
   431 => x"c048d0ff",
   432 => x"dfc278e0",
   433 => x"66cc1efa",
   434 => x"c292d44a",
   435 => x"7249e1f1",
   436 => x"eecafe81",
   437 => x"c186cc87",
   438 => x"c2c105ac",
   439 => x"4966c487",
   440 => x"1e7131c9",
   441 => x"d44a66c4",
   442 => x"e1f1c292",
   443 => x"fe817249",
   444 => x"c287dfcb",
   445 => x"c81efadf",
   446 => x"92d44a66",
   447 => x"49e1f1c2",
   448 => x"c8fe8172",
   449 => x"49d787ee",
   450 => x"87fad3ff",
   451 => x"c21ec0c8",
   452 => x"fd49fadf",
   453 => x"cc87e1e6",
   454 => x"48d0ff86",
   455 => x"f878e0c0",
   456 => x"87e7fc8e",
   457 => x"5c5b5e0e",
   458 => x"711e0e5d",
   459 => x"4cd4ff4d",
   460 => x"487e66d4",
   461 => x"06a8b7c3",
   462 => x"48c087c5",
   463 => x"7587e2c1",
   464 => x"f2d9fe49",
   465 => x"c41e7587",
   466 => x"93d44b66",
   467 => x"83e1f1c2",
   468 => x"c2fe4973",
   469 => x"83c887eb",
   470 => x"d0ff4b6b",
   471 => x"78e1c848",
   472 => x"49737cdd",
   473 => x"7199ffc3",
   474 => x"c849737c",
   475 => x"ffc329b7",
   476 => x"737c7199",
   477 => x"29b7d049",
   478 => x"7199ffc3",
   479 => x"d849737c",
   480 => x"7c7129b7",
   481 => x"7c7c7cc0",
   482 => x"7c7c7c7c",
   483 => x"7c7c7c7c",
   484 => x"78e0c07c",
   485 => x"dc1e66c4",
   486 => x"ced2ff49",
   487 => x"7386c887",
   488 => x"e4fa2648",
   489 => x"dfc21e87",
   490 => x"c149bfce",
   491 => x"d2dfc2b9",
   492 => x"48d4ff59",
   493 => x"ff78ffc3",
   494 => x"e1c048d0",
   495 => x"48d4ff78",
   496 => x"31c478c1",
   497 => x"d0ff7871",
   498 => x"78e0c048",
   499 => x"00004f26",
   500 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
