
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"dc",x"e0",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"dc",x"e0",x"c2"),
    14 => (x"48",x"d0",x"ce",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"d2",x"dc"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"c4",x"4a",x"71",x"1e"),
    47 => (x"c1",x"48",x"49",x"66"),
    48 => (x"58",x"a6",x"c8",x"88"),
    49 => (x"d6",x"02",x"99",x"71"),
    50 => (x"48",x"d4",x"ff",x"87"),
    51 => (x"68",x"78",x"ff",x"c3"),
    52 => (x"49",x"66",x"c4",x"52"),
    53 => (x"c8",x"88",x"c1",x"48"),
    54 => (x"99",x"71",x"58",x"a6"),
    55 => (x"26",x"87",x"ea",x"05"),
    56 => (x"1e",x"73",x"1e",x"4f"),
    57 => (x"c3",x"4b",x"d4",x"ff"),
    58 => (x"4a",x"6b",x"7b",x"ff"),
    59 => (x"6b",x"7b",x"ff",x"c3"),
    60 => (x"72",x"32",x"c8",x"49"),
    61 => (x"7b",x"ff",x"c3",x"b1"),
    62 => (x"31",x"c8",x"4a",x"6b"),
    63 => (x"ff",x"c3",x"b2",x"71"),
    64 => (x"c8",x"49",x"6b",x"7b"),
    65 => (x"71",x"b1",x"72",x"32"),
    66 => (x"26",x"87",x"c4",x"48"),
    67 => (x"26",x"4c",x"26",x"4d"),
    68 => (x"0e",x"4f",x"26",x"4b"),
    69 => (x"5d",x"5c",x"5b",x"5e"),
    70 => (x"ff",x"4a",x"71",x"0e"),
    71 => (x"49",x"72",x"4c",x"d4"),
    72 => (x"71",x"99",x"ff",x"c3"),
    73 => (x"d0",x"ce",x"c2",x"7c"),
    74 => (x"87",x"c8",x"05",x"bf"),
    75 => (x"c9",x"48",x"66",x"d0"),
    76 => (x"58",x"a6",x"d4",x"30"),
    77 => (x"d8",x"49",x"66",x"d0"),
    78 => (x"99",x"ff",x"c3",x"29"),
    79 => (x"66",x"d0",x"7c",x"71"),
    80 => (x"c3",x"29",x"d0",x"49"),
    81 => (x"7c",x"71",x"99",x"ff"),
    82 => (x"c8",x"49",x"66",x"d0"),
    83 => (x"99",x"ff",x"c3",x"29"),
    84 => (x"66",x"d0",x"7c",x"71"),
    85 => (x"99",x"ff",x"c3",x"49"),
    86 => (x"49",x"72",x"7c",x"71"),
    87 => (x"ff",x"c3",x"29",x"d0"),
    88 => (x"6c",x"7c",x"71",x"99"),
    89 => (x"ff",x"f0",x"c9",x"4b"),
    90 => (x"ab",x"ff",x"c3",x"4d"),
    91 => (x"c3",x"87",x"d0",x"05"),
    92 => (x"4b",x"6c",x"7c",x"ff"),
    93 => (x"c6",x"02",x"8d",x"c1"),
    94 => (x"ab",x"ff",x"c3",x"87"),
    95 => (x"73",x"87",x"f0",x"02"),
    96 => (x"87",x"c7",x"fe",x"48"),
    97 => (x"ff",x"49",x"c0",x"1e"),
    98 => (x"ff",x"c3",x"48",x"d4"),
    99 => (x"c3",x"81",x"c1",x"78"),
   100 => (x"04",x"a9",x"b7",x"c8"),
   101 => (x"4f",x"26",x"87",x"f1"),
   102 => (x"e7",x"1e",x"73",x"1e"),
   103 => (x"df",x"f8",x"c4",x"87"),
   104 => (x"c0",x"1e",x"c0",x"4b"),
   105 => (x"f7",x"c1",x"f0",x"ff"),
   106 => (x"87",x"e7",x"fd",x"49"),
   107 => (x"a8",x"c1",x"86",x"c4"),
   108 => (x"87",x"ea",x"c0",x"05"),
   109 => (x"c3",x"48",x"d4",x"ff"),
   110 => (x"c0",x"c1",x"78",x"ff"),
   111 => (x"c0",x"c0",x"c0",x"c0"),
   112 => (x"f0",x"e1",x"c0",x"1e"),
   113 => (x"fd",x"49",x"e9",x"c1"),
   114 => (x"86",x"c4",x"87",x"c9"),
   115 => (x"ca",x"05",x"98",x"70"),
   116 => (x"48",x"d4",x"ff",x"87"),
   117 => (x"c1",x"78",x"ff",x"c3"),
   118 => (x"fe",x"87",x"cb",x"48"),
   119 => (x"8b",x"c1",x"87",x"e6"),
   120 => (x"87",x"fd",x"fe",x"05"),
   121 => (x"e6",x"fc",x"48",x"c0"),
   122 => (x"1e",x"73",x"1e",x"87"),
   123 => (x"c3",x"48",x"d4",x"ff"),
   124 => (x"4b",x"d3",x"78",x"ff"),
   125 => (x"ff",x"c0",x"1e",x"c0"),
   126 => (x"49",x"c1",x"c1",x"f0"),
   127 => (x"c4",x"87",x"d4",x"fc"),
   128 => (x"05",x"98",x"70",x"86"),
   129 => (x"d4",x"ff",x"87",x"ca"),
   130 => (x"78",x"ff",x"c3",x"48"),
   131 => (x"87",x"cb",x"48",x"c1"),
   132 => (x"c1",x"87",x"f1",x"fd"),
   133 => (x"db",x"ff",x"05",x"8b"),
   134 => (x"fb",x"48",x"c0",x"87"),
   135 => (x"5e",x"0e",x"87",x"f1"),
   136 => (x"ff",x"0e",x"5c",x"5b"),
   137 => (x"db",x"fd",x"4c",x"d4"),
   138 => (x"1e",x"ea",x"c6",x"87"),
   139 => (x"c1",x"f0",x"e1",x"c0"),
   140 => (x"de",x"fb",x"49",x"c8"),
   141 => (x"c1",x"86",x"c4",x"87"),
   142 => (x"87",x"c8",x"02",x"a8"),
   143 => (x"c0",x"87",x"ea",x"fe"),
   144 => (x"87",x"e2",x"c1",x"48"),
   145 => (x"70",x"87",x"da",x"fa"),
   146 => (x"ff",x"ff",x"cf",x"49"),
   147 => (x"a9",x"ea",x"c6",x"99"),
   148 => (x"fe",x"87",x"c8",x"02"),
   149 => (x"48",x"c0",x"87",x"d3"),
   150 => (x"c3",x"87",x"cb",x"c1"),
   151 => (x"f1",x"c0",x"7c",x"ff"),
   152 => (x"87",x"f4",x"fc",x"4b"),
   153 => (x"c0",x"02",x"98",x"70"),
   154 => (x"1e",x"c0",x"87",x"eb"),
   155 => (x"c1",x"f0",x"ff",x"c0"),
   156 => (x"de",x"fa",x"49",x"fa"),
   157 => (x"70",x"86",x"c4",x"87"),
   158 => (x"87",x"d9",x"05",x"98"),
   159 => (x"6c",x"7c",x"ff",x"c3"),
   160 => (x"7c",x"ff",x"c3",x"49"),
   161 => (x"c1",x"7c",x"7c",x"7c"),
   162 => (x"c4",x"02",x"99",x"c0"),
   163 => (x"d5",x"48",x"c1",x"87"),
   164 => (x"d1",x"48",x"c0",x"87"),
   165 => (x"05",x"ab",x"c2",x"87"),
   166 => (x"48",x"c0",x"87",x"c4"),
   167 => (x"8b",x"c1",x"87",x"c8"),
   168 => (x"87",x"fd",x"fe",x"05"),
   169 => (x"e4",x"f9",x"48",x"c0"),
   170 => (x"1e",x"73",x"1e",x"87"),
   171 => (x"48",x"d0",x"ce",x"c2"),
   172 => (x"4b",x"c7",x"78",x"c1"),
   173 => (x"c2",x"48",x"d0",x"ff"),
   174 => (x"87",x"c8",x"fb",x"78"),
   175 => (x"c3",x"48",x"d0",x"ff"),
   176 => (x"c0",x"1e",x"c0",x"78"),
   177 => (x"c0",x"c1",x"d0",x"e5"),
   178 => (x"87",x"c7",x"f9",x"49"),
   179 => (x"a8",x"c1",x"86",x"c4"),
   180 => (x"4b",x"87",x"c1",x"05"),
   181 => (x"c5",x"05",x"ab",x"c2"),
   182 => (x"c0",x"48",x"c0",x"87"),
   183 => (x"8b",x"c1",x"87",x"f9"),
   184 => (x"87",x"d0",x"ff",x"05"),
   185 => (x"c2",x"87",x"f7",x"fc"),
   186 => (x"70",x"58",x"d4",x"ce"),
   187 => (x"87",x"cd",x"05",x"98"),
   188 => (x"ff",x"c0",x"1e",x"c1"),
   189 => (x"49",x"d0",x"c1",x"f0"),
   190 => (x"c4",x"87",x"d8",x"f8"),
   191 => (x"48",x"d4",x"ff",x"86"),
   192 => (x"c2",x"78",x"ff",x"c3"),
   193 => (x"ce",x"c2",x"87",x"fc"),
   194 => (x"d0",x"ff",x"58",x"d8"),
   195 => (x"ff",x"78",x"c2",x"48"),
   196 => (x"ff",x"c3",x"48",x"d4"),
   197 => (x"f7",x"48",x"c1",x"78"),
   198 => (x"5e",x"0e",x"87",x"f5"),
   199 => (x"0e",x"5d",x"5c",x"5b"),
   200 => (x"4c",x"c0",x"4b",x"71"),
   201 => (x"df",x"cd",x"ee",x"c5"),
   202 => (x"48",x"d4",x"ff",x"4a"),
   203 => (x"68",x"78",x"ff",x"c3"),
   204 => (x"a9",x"fe",x"c3",x"49"),
   205 => (x"87",x"fd",x"c0",x"05"),
   206 => (x"9b",x"73",x"4d",x"70"),
   207 => (x"d0",x"87",x"cc",x"02"),
   208 => (x"49",x"73",x"1e",x"66"),
   209 => (x"c4",x"87",x"f1",x"f5"),
   210 => (x"ff",x"87",x"d6",x"86"),
   211 => (x"d1",x"c4",x"48",x"d0"),
   212 => (x"7d",x"ff",x"c3",x"78"),
   213 => (x"c1",x"48",x"66",x"d0"),
   214 => (x"58",x"a6",x"d4",x"88"),
   215 => (x"f0",x"05",x"98",x"70"),
   216 => (x"48",x"d4",x"ff",x"87"),
   217 => (x"78",x"78",x"ff",x"c3"),
   218 => (x"c5",x"05",x"9b",x"73"),
   219 => (x"48",x"d0",x"ff",x"87"),
   220 => (x"4a",x"c1",x"78",x"d0"),
   221 => (x"05",x"8a",x"c1",x"4c"),
   222 => (x"74",x"87",x"ee",x"fe"),
   223 => (x"87",x"cb",x"f6",x"48"),
   224 => (x"71",x"1e",x"73",x"1e"),
   225 => (x"ff",x"4b",x"c0",x"4a"),
   226 => (x"ff",x"c3",x"48",x"d4"),
   227 => (x"48",x"d0",x"ff",x"78"),
   228 => (x"ff",x"78",x"c3",x"c4"),
   229 => (x"ff",x"c3",x"48",x"d4"),
   230 => (x"c0",x"1e",x"72",x"78"),
   231 => (x"d1",x"c1",x"f0",x"ff"),
   232 => (x"87",x"ef",x"f5",x"49"),
   233 => (x"98",x"70",x"86",x"c4"),
   234 => (x"c8",x"87",x"d2",x"05"),
   235 => (x"66",x"cc",x"1e",x"c0"),
   236 => (x"87",x"e6",x"fd",x"49"),
   237 => (x"4b",x"70",x"86",x"c4"),
   238 => (x"c2",x"48",x"d0",x"ff"),
   239 => (x"f5",x"48",x"73",x"78"),
   240 => (x"5e",x"0e",x"87",x"cd"),
   241 => (x"0e",x"5d",x"5c",x"5b"),
   242 => (x"ff",x"c0",x"1e",x"c0"),
   243 => (x"49",x"c9",x"c1",x"f0"),
   244 => (x"d2",x"87",x"c0",x"f5"),
   245 => (x"d8",x"ce",x"c2",x"1e"),
   246 => (x"87",x"fe",x"fc",x"49"),
   247 => (x"4c",x"c0",x"86",x"c8"),
   248 => (x"b7",x"d2",x"84",x"c1"),
   249 => (x"87",x"f8",x"04",x"ac"),
   250 => (x"97",x"d8",x"ce",x"c2"),
   251 => (x"c0",x"c3",x"49",x"bf"),
   252 => (x"a9",x"c0",x"c1",x"99"),
   253 => (x"87",x"e7",x"c0",x"05"),
   254 => (x"97",x"df",x"ce",x"c2"),
   255 => (x"31",x"d0",x"49",x"bf"),
   256 => (x"97",x"e0",x"ce",x"c2"),
   257 => (x"32",x"c8",x"4a",x"bf"),
   258 => (x"ce",x"c2",x"b1",x"72"),
   259 => (x"4a",x"bf",x"97",x"e1"),
   260 => (x"cf",x"4c",x"71",x"b1"),
   261 => (x"9c",x"ff",x"ff",x"ff"),
   262 => (x"34",x"ca",x"84",x"c1"),
   263 => (x"c2",x"87",x"e7",x"c1"),
   264 => (x"bf",x"97",x"e1",x"ce"),
   265 => (x"c6",x"31",x"c1",x"49"),
   266 => (x"e2",x"ce",x"c2",x"99"),
   267 => (x"c7",x"4a",x"bf",x"97"),
   268 => (x"b1",x"72",x"2a",x"b7"),
   269 => (x"97",x"dd",x"ce",x"c2"),
   270 => (x"cf",x"4d",x"4a",x"bf"),
   271 => (x"de",x"ce",x"c2",x"9d"),
   272 => (x"c3",x"4a",x"bf",x"97"),
   273 => (x"c2",x"32",x"ca",x"9a"),
   274 => (x"bf",x"97",x"df",x"ce"),
   275 => (x"73",x"33",x"c2",x"4b"),
   276 => (x"e0",x"ce",x"c2",x"b2"),
   277 => (x"c3",x"4b",x"bf",x"97"),
   278 => (x"b7",x"c6",x"9b",x"c0"),
   279 => (x"c2",x"b2",x"73",x"2b"),
   280 => (x"71",x"48",x"c1",x"81"),
   281 => (x"c1",x"49",x"70",x"30"),
   282 => (x"70",x"30",x"75",x"48"),
   283 => (x"c1",x"4c",x"72",x"4d"),
   284 => (x"c8",x"94",x"71",x"84"),
   285 => (x"06",x"ad",x"b7",x"c0"),
   286 => (x"34",x"c1",x"87",x"cc"),
   287 => (x"c0",x"c8",x"2d",x"b7"),
   288 => (x"ff",x"01",x"ad",x"b7"),
   289 => (x"48",x"74",x"87",x"f4"),
   290 => (x"0e",x"87",x"c0",x"f2"),
   291 => (x"5d",x"5c",x"5b",x"5e"),
   292 => (x"c2",x"86",x"f8",x"0e"),
   293 => (x"c0",x"48",x"fe",x"d6"),
   294 => (x"f6",x"ce",x"c2",x"78"),
   295 => (x"fb",x"49",x"c0",x"1e"),
   296 => (x"86",x"c4",x"87",x"de"),
   297 => (x"c5",x"05",x"98",x"70"),
   298 => (x"c9",x"48",x"c0",x"87"),
   299 => (x"4d",x"c0",x"87",x"ce"),
   300 => (x"ed",x"c0",x"7e",x"c1"),
   301 => (x"c2",x"49",x"bf",x"f3"),
   302 => (x"71",x"4a",x"ec",x"cf"),
   303 => (x"e9",x"ee",x"4b",x"c8"),
   304 => (x"05",x"98",x"70",x"87"),
   305 => (x"7e",x"c0",x"87",x"c2"),
   306 => (x"bf",x"ef",x"ed",x"c0"),
   307 => (x"c8",x"d0",x"c2",x"49"),
   308 => (x"4b",x"c8",x"71",x"4a"),
   309 => (x"70",x"87",x"d3",x"ee"),
   310 => (x"87",x"c2",x"05",x"98"),
   311 => (x"02",x"6e",x"7e",x"c0"),
   312 => (x"c2",x"87",x"fd",x"c0"),
   313 => (x"4d",x"bf",x"fc",x"d5"),
   314 => (x"9f",x"f4",x"d6",x"c2"),
   315 => (x"c5",x"48",x"7e",x"bf"),
   316 => (x"05",x"a8",x"ea",x"d6"),
   317 => (x"d5",x"c2",x"87",x"c7"),
   318 => (x"ce",x"4d",x"bf",x"fc"),
   319 => (x"ca",x"48",x"6e",x"87"),
   320 => (x"02",x"a8",x"d5",x"e9"),
   321 => (x"48",x"c0",x"87",x"c5"),
   322 => (x"c2",x"87",x"f1",x"c7"),
   323 => (x"75",x"1e",x"f6",x"ce"),
   324 => (x"87",x"ec",x"f9",x"49"),
   325 => (x"98",x"70",x"86",x"c4"),
   326 => (x"c0",x"87",x"c5",x"05"),
   327 => (x"87",x"dc",x"c7",x"48"),
   328 => (x"bf",x"ef",x"ed",x"c0"),
   329 => (x"c8",x"d0",x"c2",x"49"),
   330 => (x"4b",x"c8",x"71",x"4a"),
   331 => (x"70",x"87",x"fb",x"ec"),
   332 => (x"87",x"c8",x"05",x"98"),
   333 => (x"48",x"fe",x"d6",x"c2"),
   334 => (x"87",x"da",x"78",x"c1"),
   335 => (x"bf",x"f3",x"ed",x"c0"),
   336 => (x"ec",x"cf",x"c2",x"49"),
   337 => (x"4b",x"c8",x"71",x"4a"),
   338 => (x"70",x"87",x"df",x"ec"),
   339 => (x"c5",x"c0",x"02",x"98"),
   340 => (x"c6",x"48",x"c0",x"87"),
   341 => (x"d6",x"c2",x"87",x"e6"),
   342 => (x"49",x"bf",x"97",x"f4"),
   343 => (x"05",x"a9",x"d5",x"c1"),
   344 => (x"c2",x"87",x"cd",x"c0"),
   345 => (x"bf",x"97",x"f5",x"d6"),
   346 => (x"a9",x"ea",x"c2",x"49"),
   347 => (x"87",x"c5",x"c0",x"02"),
   348 => (x"c7",x"c6",x"48",x"c0"),
   349 => (x"f6",x"ce",x"c2",x"87"),
   350 => (x"48",x"7e",x"bf",x"97"),
   351 => (x"02",x"a8",x"e9",x"c3"),
   352 => (x"6e",x"87",x"ce",x"c0"),
   353 => (x"a8",x"eb",x"c3",x"48"),
   354 => (x"87",x"c5",x"c0",x"02"),
   355 => (x"eb",x"c5",x"48",x"c0"),
   356 => (x"c1",x"cf",x"c2",x"87"),
   357 => (x"99",x"49",x"bf",x"97"),
   358 => (x"87",x"cc",x"c0",x"05"),
   359 => (x"97",x"c2",x"cf",x"c2"),
   360 => (x"a9",x"c2",x"49",x"bf"),
   361 => (x"87",x"c5",x"c0",x"02"),
   362 => (x"cf",x"c5",x"48",x"c0"),
   363 => (x"c3",x"cf",x"c2",x"87"),
   364 => (x"c2",x"48",x"bf",x"97"),
   365 => (x"70",x"58",x"fa",x"d6"),
   366 => (x"88",x"c1",x"48",x"4c"),
   367 => (x"58",x"fe",x"d6",x"c2"),
   368 => (x"97",x"c4",x"cf",x"c2"),
   369 => (x"81",x"75",x"49",x"bf"),
   370 => (x"97",x"c5",x"cf",x"c2"),
   371 => (x"32",x"c8",x"4a",x"bf"),
   372 => (x"c2",x"7e",x"a1",x"72"),
   373 => (x"6e",x"48",x"cb",x"db"),
   374 => (x"c6",x"cf",x"c2",x"78"),
   375 => (x"c8",x"48",x"bf",x"97"),
   376 => (x"d6",x"c2",x"58",x"a6"),
   377 => (x"c2",x"02",x"bf",x"fe"),
   378 => (x"ed",x"c0",x"87",x"d4"),
   379 => (x"c2",x"49",x"bf",x"ef"),
   380 => (x"71",x"4a",x"c8",x"d0"),
   381 => (x"f1",x"e9",x"4b",x"c8"),
   382 => (x"02",x"98",x"70",x"87"),
   383 => (x"c0",x"87",x"c5",x"c0"),
   384 => (x"87",x"f8",x"c3",x"48"),
   385 => (x"bf",x"f6",x"d6",x"c2"),
   386 => (x"df",x"db",x"c2",x"4c"),
   387 => (x"db",x"cf",x"c2",x"5c"),
   388 => (x"c8",x"49",x"bf",x"97"),
   389 => (x"da",x"cf",x"c2",x"31"),
   390 => (x"a1",x"4a",x"bf",x"97"),
   391 => (x"dc",x"cf",x"c2",x"49"),
   392 => (x"d0",x"4a",x"bf",x"97"),
   393 => (x"49",x"a1",x"72",x"32"),
   394 => (x"97",x"dd",x"cf",x"c2"),
   395 => (x"32",x"d8",x"4a",x"bf"),
   396 => (x"c4",x"49",x"a1",x"72"),
   397 => (x"db",x"c2",x"91",x"66"),
   398 => (x"c2",x"81",x"bf",x"cb"),
   399 => (x"c2",x"59",x"d3",x"db"),
   400 => (x"bf",x"97",x"e3",x"cf"),
   401 => (x"c2",x"32",x"c8",x"4a"),
   402 => (x"bf",x"97",x"e2",x"cf"),
   403 => (x"c2",x"4a",x"a2",x"4b"),
   404 => (x"bf",x"97",x"e4",x"cf"),
   405 => (x"73",x"33",x"d0",x"4b"),
   406 => (x"cf",x"c2",x"4a",x"a2"),
   407 => (x"4b",x"bf",x"97",x"e5"),
   408 => (x"33",x"d8",x"9b",x"cf"),
   409 => (x"c2",x"4a",x"a2",x"73"),
   410 => (x"c2",x"5a",x"d7",x"db"),
   411 => (x"4a",x"bf",x"d3",x"db"),
   412 => (x"92",x"74",x"8a",x"c2"),
   413 => (x"48",x"d7",x"db",x"c2"),
   414 => (x"c1",x"78",x"a1",x"72"),
   415 => (x"cf",x"c2",x"87",x"ca"),
   416 => (x"49",x"bf",x"97",x"c8"),
   417 => (x"cf",x"c2",x"31",x"c8"),
   418 => (x"4a",x"bf",x"97",x"c7"),
   419 => (x"d7",x"c2",x"49",x"a1"),
   420 => (x"d7",x"c2",x"59",x"c6"),
   421 => (x"c5",x"49",x"bf",x"c2"),
   422 => (x"81",x"ff",x"c7",x"31"),
   423 => (x"db",x"c2",x"29",x"c9"),
   424 => (x"cf",x"c2",x"59",x"df"),
   425 => (x"4a",x"bf",x"97",x"cd"),
   426 => (x"cf",x"c2",x"32",x"c8"),
   427 => (x"4b",x"bf",x"97",x"cc"),
   428 => (x"66",x"c4",x"4a",x"a2"),
   429 => (x"c2",x"82",x"6e",x"92"),
   430 => (x"c2",x"5a",x"db",x"db"),
   431 => (x"c0",x"48",x"d3",x"db"),
   432 => (x"cf",x"db",x"c2",x"78"),
   433 => (x"78",x"a1",x"72",x"48"),
   434 => (x"48",x"df",x"db",x"c2"),
   435 => (x"bf",x"d3",x"db",x"c2"),
   436 => (x"e3",x"db",x"c2",x"78"),
   437 => (x"d7",x"db",x"c2",x"48"),
   438 => (x"d6",x"c2",x"78",x"bf"),
   439 => (x"c0",x"02",x"bf",x"fe"),
   440 => (x"48",x"74",x"87",x"c9"),
   441 => (x"7e",x"70",x"30",x"c4"),
   442 => (x"c2",x"87",x"c9",x"c0"),
   443 => (x"48",x"bf",x"db",x"db"),
   444 => (x"7e",x"70",x"30",x"c4"),
   445 => (x"48",x"c2",x"d7",x"c2"),
   446 => (x"48",x"c1",x"78",x"6e"),
   447 => (x"4d",x"26",x"8e",x"f8"),
   448 => (x"4b",x"26",x"4c",x"26"),
   449 => (x"5e",x"0e",x"4f",x"26"),
   450 => (x"0e",x"5d",x"5c",x"5b"),
   451 => (x"d6",x"c2",x"4a",x"71"),
   452 => (x"cb",x"02",x"bf",x"fe"),
   453 => (x"c7",x"4b",x"72",x"87"),
   454 => (x"c1",x"4c",x"72",x"2b"),
   455 => (x"87",x"c9",x"9c",x"ff"),
   456 => (x"2b",x"c8",x"4b",x"72"),
   457 => (x"ff",x"c3",x"4c",x"72"),
   458 => (x"cb",x"db",x"c2",x"9c"),
   459 => (x"ed",x"c0",x"83",x"bf"),
   460 => (x"02",x"ab",x"bf",x"eb"),
   461 => (x"ed",x"c0",x"87",x"d9"),
   462 => (x"ce",x"c2",x"5b",x"ef"),
   463 => (x"49",x"73",x"1e",x"f6"),
   464 => (x"c4",x"87",x"fd",x"f0"),
   465 => (x"05",x"98",x"70",x"86"),
   466 => (x"48",x"c0",x"87",x"c5"),
   467 => (x"c2",x"87",x"e6",x"c0"),
   468 => (x"02",x"bf",x"fe",x"d6"),
   469 => (x"49",x"74",x"87",x"d2"),
   470 => (x"ce",x"c2",x"91",x"c4"),
   471 => (x"4d",x"69",x"81",x"f6"),
   472 => (x"ff",x"ff",x"ff",x"cf"),
   473 => (x"87",x"cb",x"9d",x"ff"),
   474 => (x"91",x"c2",x"49",x"74"),
   475 => (x"81",x"f6",x"ce",x"c2"),
   476 => (x"75",x"4d",x"69",x"9f"),
   477 => (x"87",x"c6",x"fe",x"48"),
   478 => (x"5c",x"5b",x"5e",x"0e"),
   479 => (x"86",x"f8",x"0e",x"5d"),
   480 => (x"05",x"9c",x"4c",x"71"),
   481 => (x"48",x"c0",x"87",x"c5"),
   482 => (x"c8",x"87",x"c1",x"c3"),
   483 => (x"48",x"6e",x"7e",x"a4"),
   484 => (x"66",x"d8",x"78",x"c0"),
   485 => (x"d8",x"87",x"c7",x"02"),
   486 => (x"05",x"bf",x"97",x"66"),
   487 => (x"48",x"c0",x"87",x"c5"),
   488 => (x"c0",x"87",x"e9",x"c2"),
   489 => (x"c7",x"49",x"c1",x"1e"),
   490 => (x"86",x"c4",x"87",x"e6"),
   491 => (x"02",x"9d",x"4d",x"70"),
   492 => (x"c2",x"87",x"c2",x"c1"),
   493 => (x"d8",x"4a",x"c6",x"d7"),
   494 => (x"d2",x"e2",x"49",x"66"),
   495 => (x"02",x"98",x"70",x"87"),
   496 => (x"75",x"87",x"f2",x"c0"),
   497 => (x"49",x"66",x"d8",x"4a"),
   498 => (x"f7",x"e2",x"4b",x"cb"),
   499 => (x"02",x"98",x"70",x"87"),
   500 => (x"c0",x"87",x"e2",x"c0"),
   501 => (x"02",x"9d",x"75",x"1e"),
   502 => (x"a6",x"c8",x"87",x"c7"),
   503 => (x"c5",x"78",x"c0",x"48"),
   504 => (x"48",x"a6",x"c8",x"87"),
   505 => (x"66",x"c8",x"78",x"c1"),
   506 => (x"87",x"e4",x"c6",x"49"),
   507 => (x"4d",x"70",x"86",x"c4"),
   508 => (x"fe",x"fe",x"05",x"9d"),
   509 => (x"02",x"9d",x"75",x"87"),
   510 => (x"dc",x"87",x"cf",x"c1"),
   511 => (x"48",x"6e",x"49",x"a5"),
   512 => (x"a5",x"da",x"78",x"69"),
   513 => (x"48",x"a6",x"c4",x"49"),
   514 => (x"9f",x"78",x"a4",x"c4"),
   515 => (x"66",x"c4",x"48",x"69"),
   516 => (x"d6",x"c2",x"78",x"08"),
   517 => (x"d2",x"02",x"bf",x"fe"),
   518 => (x"49",x"a5",x"d4",x"87"),
   519 => (x"c0",x"49",x"69",x"9f"),
   520 => (x"71",x"99",x"ff",x"ff"),
   521 => (x"70",x"30",x"d0",x"48"),
   522 => (x"c0",x"87",x"c2",x"7e"),
   523 => (x"48",x"49",x"6e",x"7e"),
   524 => (x"80",x"bf",x"66",x"c4"),
   525 => (x"78",x"08",x"66",x"c4"),
   526 => (x"a4",x"cc",x"7c",x"c0"),
   527 => (x"bf",x"66",x"c4",x"49"),
   528 => (x"49",x"a4",x"d0",x"79"),
   529 => (x"48",x"c1",x"79",x"c0"),
   530 => (x"48",x"c0",x"87",x"c2"),
   531 => (x"ed",x"fa",x"8e",x"f8"),
   532 => (x"5b",x"5e",x"0e",x"87"),
   533 => (x"71",x"0e",x"5d",x"5c"),
   534 => (x"c1",x"02",x"9c",x"4c"),
   535 => (x"a4",x"c8",x"87",x"ca"),
   536 => (x"c1",x"02",x"69",x"49"),
   537 => (x"66",x"d0",x"87",x"c2"),
   538 => (x"82",x"49",x"6c",x"4a"),
   539 => (x"d0",x"5a",x"a6",x"d4"),
   540 => (x"c2",x"b9",x"4d",x"66"),
   541 => (x"4a",x"bf",x"fa",x"d6"),
   542 => (x"99",x"72",x"ba",x"ff"),
   543 => (x"c0",x"02",x"99",x"71"),
   544 => (x"a4",x"c4",x"87",x"e4"),
   545 => (x"f9",x"49",x"6b",x"4b"),
   546 => (x"7b",x"70",x"87",x"fc"),
   547 => (x"bf",x"f6",x"d6",x"c2"),
   548 => (x"71",x"81",x"6c",x"49"),
   549 => (x"c2",x"b9",x"75",x"7c"),
   550 => (x"4a",x"bf",x"fa",x"d6"),
   551 => (x"99",x"72",x"ba",x"ff"),
   552 => (x"ff",x"05",x"99",x"71"),
   553 => (x"7c",x"75",x"87",x"dc"),
   554 => (x"1e",x"87",x"d3",x"f9"),
   555 => (x"4b",x"71",x"1e",x"73"),
   556 => (x"87",x"c7",x"02",x"9b"),
   557 => (x"69",x"49",x"a3",x"c8"),
   558 => (x"c0",x"87",x"c5",x"05"),
   559 => (x"87",x"f7",x"c0",x"48"),
   560 => (x"bf",x"cf",x"db",x"c2"),
   561 => (x"49",x"a3",x"c4",x"4a"),
   562 => (x"89",x"c2",x"49",x"69"),
   563 => (x"bf",x"f6",x"d6",x"c2"),
   564 => (x"4a",x"a2",x"71",x"91"),
   565 => (x"bf",x"fa",x"d6",x"c2"),
   566 => (x"71",x"99",x"6b",x"49"),
   567 => (x"ed",x"c0",x"4a",x"a2"),
   568 => (x"66",x"c8",x"5a",x"ef"),
   569 => (x"ea",x"49",x"72",x"1e"),
   570 => (x"86",x"c4",x"87",x"d6"),
   571 => (x"c4",x"05",x"98",x"70"),
   572 => (x"c2",x"48",x"c0",x"87"),
   573 => (x"f8",x"48",x"c1",x"87"),
   574 => (x"73",x"1e",x"87",x"c8"),
   575 => (x"9b",x"4b",x"71",x"1e"),
   576 => (x"87",x"e4",x"c0",x"02"),
   577 => (x"5b",x"e3",x"db",x"c2"),
   578 => (x"8a",x"c2",x"4a",x"73"),
   579 => (x"bf",x"f6",x"d6",x"c2"),
   580 => (x"db",x"c2",x"92",x"49"),
   581 => (x"72",x"48",x"bf",x"cf"),
   582 => (x"e7",x"db",x"c2",x"80"),
   583 => (x"c4",x"48",x"71",x"58"),
   584 => (x"c6",x"d7",x"c2",x"30"),
   585 => (x"87",x"ed",x"c0",x"58"),
   586 => (x"48",x"df",x"db",x"c2"),
   587 => (x"bf",x"d3",x"db",x"c2"),
   588 => (x"e3",x"db",x"c2",x"78"),
   589 => (x"d7",x"db",x"c2",x"48"),
   590 => (x"d6",x"c2",x"78",x"bf"),
   591 => (x"c9",x"02",x"bf",x"fe"),
   592 => (x"f6",x"d6",x"c2",x"87"),
   593 => (x"31",x"c4",x"49",x"bf"),
   594 => (x"db",x"c2",x"87",x"c7"),
   595 => (x"c4",x"49",x"bf",x"db"),
   596 => (x"c6",x"d7",x"c2",x"31"),
   597 => (x"87",x"ea",x"f6",x"59"),
   598 => (x"5c",x"5b",x"5e",x"0e"),
   599 => (x"c0",x"4a",x"71",x"0e"),
   600 => (x"02",x"9a",x"72",x"4b"),
   601 => (x"da",x"87",x"e1",x"c0"),
   602 => (x"69",x"9f",x"49",x"a2"),
   603 => (x"fe",x"d6",x"c2",x"4b"),
   604 => (x"87",x"cf",x"02",x"bf"),
   605 => (x"9f",x"49",x"a2",x"d4"),
   606 => (x"c0",x"4c",x"49",x"69"),
   607 => (x"d0",x"9c",x"ff",x"ff"),
   608 => (x"c0",x"87",x"c2",x"34"),
   609 => (x"b3",x"49",x"74",x"4c"),
   610 => (x"ed",x"fd",x"49",x"73"),
   611 => (x"87",x"f0",x"f5",x"87"),
   612 => (x"5c",x"5b",x"5e",x"0e"),
   613 => (x"86",x"f4",x"0e",x"5d"),
   614 => (x"7e",x"c0",x"4a",x"71"),
   615 => (x"d8",x"02",x"9a",x"72"),
   616 => (x"f2",x"ce",x"c2",x"87"),
   617 => (x"c2",x"78",x"c0",x"48"),
   618 => (x"c2",x"48",x"ea",x"ce"),
   619 => (x"78",x"bf",x"e3",x"db"),
   620 => (x"48",x"ee",x"ce",x"c2"),
   621 => (x"bf",x"df",x"db",x"c2"),
   622 => (x"d3",x"d7",x"c2",x"78"),
   623 => (x"c2",x"50",x"c0",x"48"),
   624 => (x"49",x"bf",x"c2",x"d7"),
   625 => (x"bf",x"f2",x"ce",x"c2"),
   626 => (x"03",x"aa",x"71",x"4a"),
   627 => (x"72",x"87",x"c9",x"c4"),
   628 => (x"05",x"99",x"cf",x"49"),
   629 => (x"c0",x"87",x"e9",x"c0"),
   630 => (x"c2",x"48",x"eb",x"ed"),
   631 => (x"78",x"bf",x"ea",x"ce"),
   632 => (x"1e",x"f6",x"ce",x"c2"),
   633 => (x"bf",x"ea",x"ce",x"c2"),
   634 => (x"ea",x"ce",x"c2",x"49"),
   635 => (x"78",x"a1",x"c1",x"48"),
   636 => (x"87",x"cc",x"e6",x"71"),
   637 => (x"ed",x"c0",x"86",x"c4"),
   638 => (x"ce",x"c2",x"48",x"e7"),
   639 => (x"87",x"cc",x"78",x"f6"),
   640 => (x"bf",x"e7",x"ed",x"c0"),
   641 => (x"80",x"e0",x"c0",x"48"),
   642 => (x"58",x"eb",x"ed",x"c0"),
   643 => (x"bf",x"f2",x"ce",x"c2"),
   644 => (x"c2",x"80",x"c1",x"48"),
   645 => (x"27",x"58",x"f6",x"ce"),
   646 => (x"00",x"00",x"0b",x"67"),
   647 => (x"4d",x"bf",x"97",x"bf"),
   648 => (x"e3",x"c2",x"02",x"9d"),
   649 => (x"ad",x"e5",x"c3",x"87"),
   650 => (x"87",x"dc",x"c2",x"02"),
   651 => (x"bf",x"e7",x"ed",x"c0"),
   652 => (x"49",x"a3",x"cb",x"4b"),
   653 => (x"ac",x"cf",x"4c",x"11"),
   654 => (x"87",x"d2",x"c1",x"05"),
   655 => (x"99",x"df",x"49",x"75"),
   656 => (x"91",x"cd",x"89",x"c1"),
   657 => (x"81",x"c6",x"d7",x"c2"),
   658 => (x"12",x"4a",x"a3",x"c1"),
   659 => (x"4a",x"a3",x"c3",x"51"),
   660 => (x"a3",x"c5",x"51",x"12"),
   661 => (x"c7",x"51",x"12",x"4a"),
   662 => (x"51",x"12",x"4a",x"a3"),
   663 => (x"12",x"4a",x"a3",x"c9"),
   664 => (x"4a",x"a3",x"ce",x"51"),
   665 => (x"a3",x"d0",x"51",x"12"),
   666 => (x"d2",x"51",x"12",x"4a"),
   667 => (x"51",x"12",x"4a",x"a3"),
   668 => (x"12",x"4a",x"a3",x"d4"),
   669 => (x"4a",x"a3",x"d6",x"51"),
   670 => (x"a3",x"d8",x"51",x"12"),
   671 => (x"dc",x"51",x"12",x"4a"),
   672 => (x"51",x"12",x"4a",x"a3"),
   673 => (x"12",x"4a",x"a3",x"de"),
   674 => (x"c0",x"7e",x"c1",x"51"),
   675 => (x"49",x"74",x"87",x"fa"),
   676 => (x"c0",x"05",x"99",x"c8"),
   677 => (x"49",x"74",x"87",x"eb"),
   678 => (x"d1",x"05",x"99",x"d0"),
   679 => (x"02",x"66",x"dc",x"87"),
   680 => (x"73",x"87",x"cb",x"c0"),
   681 => (x"0f",x"66",x"dc",x"49"),
   682 => (x"c0",x"02",x"98",x"70"),
   683 => (x"05",x"6e",x"87",x"d3"),
   684 => (x"c2",x"87",x"c6",x"c0"),
   685 => (x"c0",x"48",x"c6",x"d7"),
   686 => (x"e7",x"ed",x"c0",x"50"),
   687 => (x"e1",x"c2",x"48",x"bf"),
   688 => (x"d3",x"d7",x"c2",x"87"),
   689 => (x"7e",x"50",x"c0",x"48"),
   690 => (x"bf",x"c2",x"d7",x"c2"),
   691 => (x"f2",x"ce",x"c2",x"49"),
   692 => (x"aa",x"71",x"4a",x"bf"),
   693 => (x"87",x"f7",x"fb",x"04"),
   694 => (x"bf",x"e3",x"db",x"c2"),
   695 => (x"87",x"c8",x"c0",x"05"),
   696 => (x"bf",x"fe",x"d6",x"c2"),
   697 => (x"87",x"f8",x"c1",x"02"),
   698 => (x"bf",x"ee",x"ce",x"c2"),
   699 => (x"87",x"d6",x"f0",x"49"),
   700 => (x"ce",x"c2",x"49",x"70"),
   701 => (x"a6",x"c4",x"59",x"f2"),
   702 => (x"ee",x"ce",x"c2",x"48"),
   703 => (x"d6",x"c2",x"78",x"bf"),
   704 => (x"c0",x"02",x"bf",x"fe"),
   705 => (x"66",x"c4",x"87",x"d8"),
   706 => (x"ff",x"ff",x"cf",x"49"),
   707 => (x"a9",x"99",x"f8",x"ff"),
   708 => (x"87",x"c5",x"c0",x"02"),
   709 => (x"e1",x"c0",x"4c",x"c0"),
   710 => (x"c0",x"4c",x"c1",x"87"),
   711 => (x"66",x"c4",x"87",x"dc"),
   712 => (x"f8",x"ff",x"cf",x"49"),
   713 => (x"c0",x"02",x"a9",x"99"),
   714 => (x"a6",x"c8",x"87",x"c8"),
   715 => (x"c0",x"78",x"c0",x"48"),
   716 => (x"a6",x"c8",x"87",x"c5"),
   717 => (x"c8",x"78",x"c1",x"48"),
   718 => (x"9c",x"74",x"4c",x"66"),
   719 => (x"87",x"e0",x"c0",x"05"),
   720 => (x"c2",x"49",x"66",x"c4"),
   721 => (x"f6",x"d6",x"c2",x"89"),
   722 => (x"c2",x"91",x"4a",x"bf"),
   723 => (x"4a",x"bf",x"cf",x"db"),
   724 => (x"48",x"ea",x"ce",x"c2"),
   725 => (x"c2",x"78",x"a1",x"72"),
   726 => (x"c0",x"48",x"f2",x"ce"),
   727 => (x"87",x"df",x"f9",x"78"),
   728 => (x"8e",x"f4",x"48",x"c0"),
   729 => (x"00",x"87",x"d7",x"ee"),
   730 => (x"ff",x"00",x"00",x"00"),
   731 => (x"77",x"ff",x"ff",x"ff"),
   732 => (x"80",x"00",x"00",x"0b"),
   733 => (x"46",x"00",x"00",x"0b"),
   734 => (x"32",x"33",x"54",x"41"),
   735 => (x"00",x"20",x"20",x"20"),
   736 => (x"31",x"54",x"41",x"46"),
   737 => (x"20",x"20",x"20",x"36"),
   738 => (x"d4",x"ff",x"1e",x"00"),
   739 => (x"78",x"ff",x"c3",x"48"),
   740 => (x"4f",x"26",x"48",x"68"),
   741 => (x"48",x"d4",x"ff",x"1e"),
   742 => (x"ff",x"78",x"ff",x"c3"),
   743 => (x"e1",x"c0",x"48",x"d0"),
   744 => (x"48",x"d4",x"ff",x"78"),
   745 => (x"db",x"c2",x"78",x"d4"),
   746 => (x"d4",x"ff",x"48",x"e7"),
   747 => (x"4f",x"26",x"50",x"bf"),
   748 => (x"48",x"d0",x"ff",x"1e"),
   749 => (x"26",x"78",x"e0",x"c0"),
   750 => (x"cc",x"ff",x"1e",x"4f"),
   751 => (x"99",x"49",x"70",x"87"),
   752 => (x"c0",x"87",x"c6",x"02"),
   753 => (x"f1",x"05",x"a9",x"fb"),
   754 => (x"26",x"48",x"71",x"87"),
   755 => (x"5b",x"5e",x"0e",x"4f"),
   756 => (x"4b",x"71",x"0e",x"5c"),
   757 => (x"f0",x"fe",x"4c",x"c0"),
   758 => (x"99",x"49",x"70",x"87"),
   759 => (x"87",x"f9",x"c0",x"02"),
   760 => (x"02",x"a9",x"ec",x"c0"),
   761 => (x"c0",x"87",x"f2",x"c0"),
   762 => (x"c0",x"02",x"a9",x"fb"),
   763 => (x"66",x"cc",x"87",x"eb"),
   764 => (x"c7",x"03",x"ac",x"b7"),
   765 => (x"02",x"66",x"d0",x"87"),
   766 => (x"53",x"71",x"87",x"c2"),
   767 => (x"c2",x"02",x"99",x"71"),
   768 => (x"fe",x"84",x"c1",x"87"),
   769 => (x"49",x"70",x"87",x"c3"),
   770 => (x"87",x"cd",x"02",x"99"),
   771 => (x"02",x"a9",x"ec",x"c0"),
   772 => (x"fb",x"c0",x"87",x"c7"),
   773 => (x"d5",x"ff",x"05",x"a9"),
   774 => (x"02",x"66",x"d0",x"87"),
   775 => (x"97",x"c0",x"87",x"c3"),
   776 => (x"a9",x"ec",x"c0",x"7b"),
   777 => (x"74",x"87",x"c4",x"05"),
   778 => (x"74",x"87",x"c5",x"4a"),
   779 => (x"8a",x"0a",x"c0",x"4a"),
   780 => (x"87",x"c2",x"48",x"72"),
   781 => (x"4c",x"26",x"4d",x"26"),
   782 => (x"4f",x"26",x"4b",x"26"),
   783 => (x"87",x"c9",x"fd",x"1e"),
   784 => (x"c0",x"4a",x"49",x"70"),
   785 => (x"c9",x"04",x"aa",x"f0"),
   786 => (x"aa",x"f9",x"c0",x"87"),
   787 => (x"c0",x"87",x"c3",x"01"),
   788 => (x"c1",x"c1",x"8a",x"f0"),
   789 => (x"87",x"c9",x"04",x"aa"),
   790 => (x"01",x"aa",x"da",x"c1"),
   791 => (x"f7",x"c0",x"87",x"c3"),
   792 => (x"26",x"48",x"72",x"8a"),
   793 => (x"5b",x"5e",x"0e",x"4f"),
   794 => (x"4a",x"71",x"0e",x"5c"),
   795 => (x"72",x"4c",x"d4",x"ff"),
   796 => (x"87",x"e9",x"c0",x"49"),
   797 => (x"02",x"9b",x"4b",x"70"),
   798 => (x"8b",x"c1",x"87",x"c2"),
   799 => (x"c5",x"48",x"d0",x"ff"),
   800 => (x"7c",x"d5",x"c1",x"78"),
   801 => (x"31",x"c6",x"49",x"73"),
   802 => (x"97",x"f3",x"dd",x"c1"),
   803 => (x"71",x"48",x"4a",x"bf"),
   804 => (x"ff",x"7c",x"70",x"b0"),
   805 => (x"78",x"c4",x"48",x"d0"),
   806 => (x"d9",x"fe",x"48",x"73"),
   807 => (x"5b",x"5e",x"0e",x"87"),
   808 => (x"f8",x"0e",x"5d",x"5c"),
   809 => (x"c0",x"4c",x"71",x"86"),
   810 => (x"87",x"e8",x"fb",x"7e"),
   811 => (x"f5",x"c0",x"4b",x"c0"),
   812 => (x"49",x"bf",x"97",x"ca"),
   813 => (x"cf",x"04",x"a9",x"c0"),
   814 => (x"87",x"fd",x"fb",x"87"),
   815 => (x"f5",x"c0",x"83",x"c1"),
   816 => (x"49",x"bf",x"97",x"ca"),
   817 => (x"87",x"f1",x"06",x"ab"),
   818 => (x"97",x"ca",x"f5",x"c0"),
   819 => (x"87",x"cf",x"02",x"bf"),
   820 => (x"70",x"87",x"f6",x"fa"),
   821 => (x"c6",x"02",x"99",x"49"),
   822 => (x"a9",x"ec",x"c0",x"87"),
   823 => (x"c0",x"87",x"f1",x"05"),
   824 => (x"87",x"e5",x"fa",x"4b"),
   825 => (x"e0",x"fa",x"4d",x"70"),
   826 => (x"58",x"a6",x"c8",x"87"),
   827 => (x"70",x"87",x"da",x"fa"),
   828 => (x"c8",x"83",x"c1",x"4a"),
   829 => (x"69",x"97",x"49",x"a4"),
   830 => (x"c7",x"02",x"ad",x"49"),
   831 => (x"ad",x"ff",x"c0",x"87"),
   832 => (x"87",x"e7",x"c0",x"05"),
   833 => (x"97",x"49",x"a4",x"c9"),
   834 => (x"66",x"c4",x"49",x"69"),
   835 => (x"87",x"c7",x"02",x"a9"),
   836 => (x"a8",x"ff",x"c0",x"48"),
   837 => (x"ca",x"87",x"d4",x"05"),
   838 => (x"69",x"97",x"49",x"a4"),
   839 => (x"c6",x"02",x"aa",x"49"),
   840 => (x"aa",x"ff",x"c0",x"87"),
   841 => (x"c1",x"87",x"c4",x"05"),
   842 => (x"c0",x"87",x"d0",x"7e"),
   843 => (x"c6",x"02",x"ad",x"ec"),
   844 => (x"ad",x"fb",x"c0",x"87"),
   845 => (x"c0",x"87",x"c4",x"05"),
   846 => (x"6e",x"7e",x"c1",x"4b"),
   847 => (x"87",x"e1",x"fe",x"02"),
   848 => (x"73",x"87",x"ed",x"f9"),
   849 => (x"fb",x"8e",x"f8",x"48"),
   850 => (x"0e",x"00",x"87",x"ea"),
   851 => (x"5d",x"5c",x"5b",x"5e"),
   852 => (x"71",x"86",x"f8",x"0e"),
   853 => (x"4b",x"d4",x"ff",x"4d"),
   854 => (x"db",x"c2",x"1e",x"75"),
   855 => (x"d7",x"e8",x"49",x"ec"),
   856 => (x"70",x"86",x"c4",x"87"),
   857 => (x"cc",x"c4",x"02",x"98"),
   858 => (x"48",x"a6",x"c4",x"87"),
   859 => (x"bf",x"f5",x"dd",x"c1"),
   860 => (x"fb",x"49",x"75",x"78"),
   861 => (x"d0",x"ff",x"87",x"ef"),
   862 => (x"c1",x"78",x"c5",x"48"),
   863 => (x"4a",x"c0",x"7b",x"d6"),
   864 => (x"11",x"49",x"a2",x"75"),
   865 => (x"cb",x"82",x"c1",x"7b"),
   866 => (x"f3",x"04",x"aa",x"b7"),
   867 => (x"c3",x"4a",x"cc",x"87"),
   868 => (x"82",x"c1",x"7b",x"ff"),
   869 => (x"aa",x"b7",x"e0",x"c0"),
   870 => (x"ff",x"87",x"f4",x"04"),
   871 => (x"78",x"c4",x"48",x"d0"),
   872 => (x"c5",x"7b",x"ff",x"c3"),
   873 => (x"7b",x"d3",x"c1",x"78"),
   874 => (x"78",x"c4",x"7b",x"c1"),
   875 => (x"b7",x"c0",x"48",x"66"),
   876 => (x"f0",x"c2",x"06",x"a8"),
   877 => (x"f4",x"db",x"c2",x"87"),
   878 => (x"66",x"c4",x"4c",x"bf"),
   879 => (x"c8",x"88",x"74",x"48"),
   880 => (x"9c",x"74",x"58",x"a6"),
   881 => (x"87",x"f9",x"c1",x"02"),
   882 => (x"7e",x"f6",x"ce",x"c2"),
   883 => (x"8c",x"4d",x"c0",x"c8"),
   884 => (x"03",x"ac",x"b7",x"c0"),
   885 => (x"c0",x"c8",x"87",x"c6"),
   886 => (x"4c",x"c0",x"4d",x"a4"),
   887 => (x"97",x"e7",x"db",x"c2"),
   888 => (x"99",x"d0",x"49",x"bf"),
   889 => (x"c0",x"87",x"d1",x"02"),
   890 => (x"ec",x"db",x"c2",x"1e"),
   891 => (x"87",x"fb",x"ea",x"49"),
   892 => (x"49",x"70",x"86",x"c4"),
   893 => (x"87",x"ee",x"c0",x"4a"),
   894 => (x"1e",x"f6",x"ce",x"c2"),
   895 => (x"49",x"ec",x"db",x"c2"),
   896 => (x"c4",x"87",x"e8",x"ea"),
   897 => (x"4a",x"49",x"70",x"86"),
   898 => (x"c8",x"48",x"d0",x"ff"),
   899 => (x"d4",x"c1",x"78",x"c5"),
   900 => (x"bf",x"97",x"6e",x"7b"),
   901 => (x"c1",x"48",x"6e",x"7b"),
   902 => (x"c1",x"7e",x"70",x"80"),
   903 => (x"f0",x"ff",x"05",x"8d"),
   904 => (x"48",x"d0",x"ff",x"87"),
   905 => (x"9a",x"72",x"78",x"c4"),
   906 => (x"c0",x"87",x"c5",x"05"),
   907 => (x"87",x"c7",x"c1",x"48"),
   908 => (x"db",x"c2",x"1e",x"c1"),
   909 => (x"d8",x"e8",x"49",x"ec"),
   910 => (x"74",x"86",x"c4",x"87"),
   911 => (x"c7",x"fe",x"05",x"9c"),
   912 => (x"48",x"66",x"c4",x"87"),
   913 => (x"06",x"a8",x"b7",x"c0"),
   914 => (x"db",x"c2",x"87",x"d1"),
   915 => (x"78",x"c0",x"48",x"ec"),
   916 => (x"78",x"c0",x"80",x"d0"),
   917 => (x"db",x"c2",x"80",x"f4"),
   918 => (x"c4",x"78",x"bf",x"f8"),
   919 => (x"b7",x"c0",x"48",x"66"),
   920 => (x"d0",x"fd",x"01",x"a8"),
   921 => (x"48",x"d0",x"ff",x"87"),
   922 => (x"d3",x"c1",x"78",x"c5"),
   923 => (x"c4",x"7b",x"c0",x"7b"),
   924 => (x"c2",x"48",x"c1",x"78"),
   925 => (x"f8",x"48",x"c0",x"87"),
   926 => (x"26",x"4d",x"26",x"8e"),
   927 => (x"26",x"4b",x"26",x"4c"),
   928 => (x"5b",x"5e",x"0e",x"4f"),
   929 => (x"1e",x"0e",x"5d",x"5c"),
   930 => (x"4c",x"c0",x"4b",x"71"),
   931 => (x"c0",x"04",x"ab",x"4d"),
   932 => (x"f2",x"c0",x"87",x"e8"),
   933 => (x"9d",x"75",x"1e",x"dd"),
   934 => (x"c0",x"87",x"c4",x"02"),
   935 => (x"c1",x"87",x"c2",x"4a"),
   936 => (x"eb",x"49",x"72",x"4a"),
   937 => (x"86",x"c4",x"87",x"ea"),
   938 => (x"84",x"c1",x"7e",x"70"),
   939 => (x"87",x"c2",x"05",x"6e"),
   940 => (x"85",x"c1",x"4c",x"73"),
   941 => (x"ff",x"06",x"ac",x"73"),
   942 => (x"48",x"6e",x"87",x"d8"),
   943 => (x"87",x"f9",x"fe",x"26"),
   944 => (x"c4",x"4a",x"71",x"1e"),
   945 => (x"87",x"c5",x"05",x"66"),
   946 => (x"fe",x"f9",x"49",x"72"),
   947 => (x"0e",x"4f",x"26",x"87"),
   948 => (x"5d",x"5c",x"5b",x"5e"),
   949 => (x"4c",x"71",x"1e",x"0e"),
   950 => (x"c2",x"91",x"de",x"49"),
   951 => (x"71",x"4d",x"d4",x"dc"),
   952 => (x"02",x"6d",x"97",x"85"),
   953 => (x"c2",x"87",x"dc",x"c1"),
   954 => (x"4a",x"bf",x"c0",x"dc"),
   955 => (x"49",x"72",x"82",x"74"),
   956 => (x"70",x"87",x"ce",x"fe"),
   957 => (x"c0",x"02",x"6e",x"7e"),
   958 => (x"dc",x"c2",x"87",x"f2"),
   959 => (x"4a",x"6e",x"4b",x"c8"),
   960 => (x"c6",x"ff",x"49",x"cb"),
   961 => (x"4b",x"74",x"87",x"e2"),
   962 => (x"de",x"c1",x"93",x"cb"),
   963 => (x"83",x"c4",x"83",x"c7"),
   964 => (x"7b",x"c7",x"fd",x"c0"),
   965 => (x"c1",x"c1",x"49",x"74"),
   966 => (x"7b",x"75",x"87",x"e7"),
   967 => (x"97",x"f4",x"dd",x"c1"),
   968 => (x"c2",x"1e",x"49",x"bf"),
   969 => (x"fe",x"49",x"c8",x"dc"),
   970 => (x"86",x"c4",x"87",x"d6"),
   971 => (x"c1",x"c1",x"49",x"74"),
   972 => (x"49",x"c0",x"87",x"cf"),
   973 => (x"87",x"ee",x"c2",x"c1"),
   974 => (x"48",x"e8",x"db",x"c2"),
   975 => (x"49",x"c1",x"78",x"c0"),
   976 => (x"26",x"87",x"d9",x"dd"),
   977 => (x"4c",x"87",x"f2",x"fc"),
   978 => (x"69",x"64",x"61",x"6f"),
   979 => (x"2e",x"2e",x"67",x"6e"),
   980 => (x"5e",x"0e",x"00",x"2e"),
   981 => (x"71",x"0e",x"5c",x"5b"),
   982 => (x"dc",x"c2",x"4a",x"4b"),
   983 => (x"72",x"82",x"bf",x"c0"),
   984 => (x"87",x"dd",x"fc",x"49"),
   985 => (x"02",x"9c",x"4c",x"70"),
   986 => (x"e7",x"49",x"87",x"c4"),
   987 => (x"dc",x"c2",x"87",x"ea"),
   988 => (x"78",x"c0",x"48",x"c0"),
   989 => (x"e3",x"dc",x"49",x"c1"),
   990 => (x"87",x"ff",x"fb",x"87"),
   991 => (x"5c",x"5b",x"5e",x"0e"),
   992 => (x"86",x"f4",x"0e",x"5d"),
   993 => (x"4d",x"f6",x"ce",x"c2"),
   994 => (x"a6",x"c4",x"4c",x"c0"),
   995 => (x"c2",x"78",x"c0",x"48"),
   996 => (x"49",x"bf",x"c0",x"dc"),
   997 => (x"c1",x"06",x"a9",x"c0"),
   998 => (x"ce",x"c2",x"87",x"c1"),
   999 => (x"02",x"98",x"48",x"f6"),
  1000 => (x"c0",x"87",x"f8",x"c0"),
  1001 => (x"c8",x"1e",x"dd",x"f2"),
  1002 => (x"87",x"c7",x"02",x"66"),
  1003 => (x"c0",x"48",x"a6",x"c4"),
  1004 => (x"c4",x"87",x"c5",x"78"),
  1005 => (x"78",x"c1",x"48",x"a6"),
  1006 => (x"e7",x"49",x"66",x"c4"),
  1007 => (x"86",x"c4",x"87",x"d2"),
  1008 => (x"84",x"c1",x"4d",x"70"),
  1009 => (x"c1",x"48",x"66",x"c4"),
  1010 => (x"58",x"a6",x"c8",x"80"),
  1011 => (x"bf",x"c0",x"dc",x"c2"),
  1012 => (x"c6",x"03",x"ac",x"49"),
  1013 => (x"05",x"9d",x"75",x"87"),
  1014 => (x"c0",x"87",x"c8",x"ff"),
  1015 => (x"02",x"9d",x"75",x"4c"),
  1016 => (x"c0",x"87",x"e0",x"c3"),
  1017 => (x"c8",x"1e",x"dd",x"f2"),
  1018 => (x"87",x"c7",x"02",x"66"),
  1019 => (x"c0",x"48",x"a6",x"cc"),
  1020 => (x"cc",x"87",x"c5",x"78"),
  1021 => (x"78",x"c1",x"48",x"a6"),
  1022 => (x"e6",x"49",x"66",x"cc"),
  1023 => (x"86",x"c4",x"87",x"d2"),
  1024 => (x"02",x"6e",x"7e",x"70"),
  1025 => (x"6e",x"87",x"e9",x"c2"),
  1026 => (x"97",x"81",x"cb",x"49"),
  1027 => (x"99",x"d0",x"49",x"69"),
  1028 => (x"87",x"d6",x"c1",x"02"),
  1029 => (x"4a",x"d2",x"fd",x"c0"),
  1030 => (x"91",x"cb",x"49",x"74"),
  1031 => (x"81",x"c7",x"de",x"c1"),
  1032 => (x"81",x"c8",x"79",x"72"),
  1033 => (x"74",x"51",x"ff",x"c3"),
  1034 => (x"c2",x"91",x"de",x"49"),
  1035 => (x"71",x"4d",x"d4",x"dc"),
  1036 => (x"97",x"c1",x"c2",x"85"),
  1037 => (x"49",x"a5",x"c1",x"7d"),
  1038 => (x"c2",x"51",x"e0",x"c0"),
  1039 => (x"bf",x"97",x"c6",x"d7"),
  1040 => (x"c1",x"87",x"d2",x"02"),
  1041 => (x"4b",x"a5",x"c2",x"84"),
  1042 => (x"4a",x"c6",x"d7",x"c2"),
  1043 => (x"c1",x"ff",x"49",x"db"),
  1044 => (x"db",x"c1",x"87",x"d6"),
  1045 => (x"49",x"a5",x"cd",x"87"),
  1046 => (x"84",x"c1",x"51",x"c0"),
  1047 => (x"6e",x"4b",x"a5",x"c2"),
  1048 => (x"ff",x"49",x"cb",x"4a"),
  1049 => (x"c1",x"87",x"c1",x"c1"),
  1050 => (x"fb",x"c0",x"87",x"c6"),
  1051 => (x"49",x"74",x"4a",x"cf"),
  1052 => (x"de",x"c1",x"91",x"cb"),
  1053 => (x"79",x"72",x"81",x"c7"),
  1054 => (x"97",x"c6",x"d7",x"c2"),
  1055 => (x"87",x"d8",x"02",x"bf"),
  1056 => (x"91",x"de",x"49",x"74"),
  1057 => (x"dc",x"c2",x"84",x"c1"),
  1058 => (x"83",x"71",x"4b",x"d4"),
  1059 => (x"4a",x"c6",x"d7",x"c2"),
  1060 => (x"c0",x"ff",x"49",x"dd"),
  1061 => (x"87",x"d8",x"87",x"d2"),
  1062 => (x"93",x"de",x"4b",x"74"),
  1063 => (x"83",x"d4",x"dc",x"c2"),
  1064 => (x"c0",x"49",x"a3",x"cb"),
  1065 => (x"73",x"84",x"c1",x"51"),
  1066 => (x"49",x"cb",x"4a",x"6e"),
  1067 => (x"87",x"f8",x"ff",x"fe"),
  1068 => (x"c1",x"48",x"66",x"c4"),
  1069 => (x"58",x"a6",x"c8",x"80"),
  1070 => (x"c0",x"03",x"ac",x"c7"),
  1071 => (x"05",x"6e",x"87",x"c5"),
  1072 => (x"74",x"87",x"e0",x"fc"),
  1073 => (x"f6",x"8e",x"f4",x"48"),
  1074 => (x"73",x"1e",x"87",x"ef"),
  1075 => (x"49",x"4b",x"71",x"1e"),
  1076 => (x"de",x"c1",x"91",x"cb"),
  1077 => (x"a1",x"c8",x"81",x"c7"),
  1078 => (x"f3",x"dd",x"c1",x"4a"),
  1079 => (x"c9",x"50",x"12",x"48"),
  1080 => (x"f5",x"c0",x"4a",x"a1"),
  1081 => (x"50",x"12",x"48",x"ca"),
  1082 => (x"dd",x"c1",x"81",x"ca"),
  1083 => (x"50",x"11",x"48",x"f4"),
  1084 => (x"97",x"f4",x"dd",x"c1"),
  1085 => (x"c0",x"1e",x"49",x"bf"),
  1086 => (x"87",x"c4",x"f7",x"49"),
  1087 => (x"48",x"e8",x"db",x"c2"),
  1088 => (x"49",x"c1",x"78",x"de"),
  1089 => (x"26",x"87",x"d5",x"d6"),
  1090 => (x"1e",x"87",x"f2",x"f5"),
  1091 => (x"cb",x"49",x"4a",x"71"),
  1092 => (x"c7",x"de",x"c1",x"91"),
  1093 => (x"11",x"81",x"c8",x"81"),
  1094 => (x"ec",x"db",x"c2",x"48"),
  1095 => (x"c0",x"dc",x"c2",x"58"),
  1096 => (x"c1",x"78",x"c0",x"48"),
  1097 => (x"87",x"f4",x"d5",x"49"),
  1098 => (x"c0",x"1e",x"4f",x"26"),
  1099 => (x"f5",x"fa",x"c0",x"49"),
  1100 => (x"1e",x"4f",x"26",x"87"),
  1101 => (x"d2",x"02",x"99",x"71"),
  1102 => (x"dc",x"df",x"c1",x"87"),
  1103 => (x"f7",x"50",x"c0",x"48"),
  1104 => (x"cb",x"c4",x"c1",x"80"),
  1105 => (x"c0",x"de",x"c1",x"40"),
  1106 => (x"c1",x"87",x"ce",x"78"),
  1107 => (x"c1",x"48",x"d8",x"df"),
  1108 => (x"fc",x"78",x"f9",x"dd"),
  1109 => (x"ea",x"c4",x"c1",x"80"),
  1110 => (x"0e",x"4f",x"26",x"78"),
  1111 => (x"0e",x"5c",x"5b",x"5e"),
  1112 => (x"cb",x"4a",x"4c",x"71"),
  1113 => (x"c7",x"de",x"c1",x"92"),
  1114 => (x"49",x"a2",x"c8",x"82"),
  1115 => (x"97",x"4b",x"a2",x"c9"),
  1116 => (x"97",x"1e",x"4b",x"6b"),
  1117 => (x"ca",x"1e",x"49",x"69"),
  1118 => (x"c0",x"49",x"12",x"82"),
  1119 => (x"c0",x"87",x"f0",x"e5"),
  1120 => (x"87",x"d8",x"d4",x"49"),
  1121 => (x"f7",x"c0",x"49",x"74"),
  1122 => (x"8e",x"f8",x"87",x"f7"),
  1123 => (x"1e",x"87",x"ec",x"f3"),
  1124 => (x"4b",x"71",x"1e",x"73"),
  1125 => (x"87",x"c3",x"ff",x"49"),
  1126 => (x"fe",x"fe",x"49",x"73"),
  1127 => (x"87",x"dd",x"f3",x"87"),
  1128 => (x"71",x"1e",x"73",x"1e"),
  1129 => (x"4a",x"a3",x"c6",x"4b"),
  1130 => (x"c1",x"87",x"db",x"02"),
  1131 => (x"87",x"d6",x"02",x"8a"),
  1132 => (x"da",x"c1",x"02",x"8a"),
  1133 => (x"c0",x"02",x"8a",x"87"),
  1134 => (x"02",x"8a",x"87",x"fc"),
  1135 => (x"8a",x"87",x"e1",x"c0"),
  1136 => (x"c1",x"87",x"cb",x"02"),
  1137 => (x"49",x"c7",x"87",x"db"),
  1138 => (x"c1",x"87",x"c0",x"fd"),
  1139 => (x"dc",x"c2",x"87",x"de"),
  1140 => (x"c1",x"02",x"bf",x"c0"),
  1141 => (x"c1",x"48",x"87",x"cb"),
  1142 => (x"c4",x"dc",x"c2",x"88"),
  1143 => (x"87",x"c1",x"c1",x"58"),
  1144 => (x"bf",x"c4",x"dc",x"c2"),
  1145 => (x"87",x"f9",x"c0",x"02"),
  1146 => (x"bf",x"c0",x"dc",x"c2"),
  1147 => (x"c2",x"80",x"c1",x"48"),
  1148 => (x"c0",x"58",x"c4",x"dc"),
  1149 => (x"dc",x"c2",x"87",x"eb"),
  1150 => (x"c6",x"49",x"bf",x"c0"),
  1151 => (x"c4",x"dc",x"c2",x"89"),
  1152 => (x"a9",x"b7",x"c0",x"59"),
  1153 => (x"c2",x"87",x"da",x"03"),
  1154 => (x"c0",x"48",x"c0",x"dc"),
  1155 => (x"c2",x"87",x"d2",x"78"),
  1156 => (x"02",x"bf",x"c4",x"dc"),
  1157 => (x"dc",x"c2",x"87",x"cb"),
  1158 => (x"c6",x"48",x"bf",x"c0"),
  1159 => (x"c4",x"dc",x"c2",x"80"),
  1160 => (x"d1",x"49",x"c0",x"58"),
  1161 => (x"49",x"73",x"87",x"f6"),
  1162 => (x"87",x"d5",x"f5",x"c0"),
  1163 => (x"0e",x"87",x"ce",x"f1"),
  1164 => (x"5d",x"5c",x"5b",x"5e"),
  1165 => (x"86",x"d0",x"ff",x"0e"),
  1166 => (x"c8",x"59",x"a6",x"dc"),
  1167 => (x"78",x"c0",x"48",x"a6"),
  1168 => (x"c4",x"c1",x"80",x"c4"),
  1169 => (x"80",x"c4",x"78",x"66"),
  1170 => (x"80",x"c4",x"78",x"c1"),
  1171 => (x"dc",x"c2",x"78",x"c1"),
  1172 => (x"78",x"c1",x"48",x"c4"),
  1173 => (x"bf",x"e8",x"db",x"c2"),
  1174 => (x"05",x"a8",x"de",x"48"),
  1175 => (x"db",x"f4",x"87",x"cb"),
  1176 => (x"cc",x"49",x"70",x"87"),
  1177 => (x"f2",x"cf",x"59",x"a6"),
  1178 => (x"87",x"e8",x"e4",x"87"),
  1179 => (x"e4",x"87",x"ca",x"e5"),
  1180 => (x"4c",x"70",x"87",x"d7"),
  1181 => (x"02",x"ac",x"fb",x"c0"),
  1182 => (x"d8",x"87",x"fb",x"c1"),
  1183 => (x"ed",x"c1",x"05",x"66"),
  1184 => (x"66",x"c0",x"c1",x"87"),
  1185 => (x"6a",x"82",x"c4",x"4a"),
  1186 => (x"c1",x"1e",x"72",x"7e"),
  1187 => (x"c4",x"48",x"d0",x"da"),
  1188 => (x"a1",x"c8",x"49",x"66"),
  1189 => (x"71",x"41",x"20",x"4a"),
  1190 => (x"87",x"f9",x"05",x"aa"),
  1191 => (x"4a",x"26",x"51",x"10"),
  1192 => (x"48",x"66",x"c0",x"c1"),
  1193 => (x"78",x"ca",x"c3",x"c1"),
  1194 => (x"81",x"c7",x"49",x"6a"),
  1195 => (x"c0",x"c1",x"51",x"74"),
  1196 => (x"81",x"c8",x"49",x"66"),
  1197 => (x"c0",x"c1",x"51",x"c1"),
  1198 => (x"81",x"c9",x"49",x"66"),
  1199 => (x"c0",x"c1",x"51",x"c0"),
  1200 => (x"81",x"ca",x"49",x"66"),
  1201 => (x"1e",x"c1",x"51",x"c0"),
  1202 => (x"49",x"6a",x"1e",x"d8"),
  1203 => (x"fc",x"e3",x"81",x"c8"),
  1204 => (x"c1",x"86",x"c8",x"87"),
  1205 => (x"c0",x"48",x"66",x"c4"),
  1206 => (x"87",x"c7",x"01",x"a8"),
  1207 => (x"c1",x"48",x"a6",x"c8"),
  1208 => (x"c1",x"87",x"ce",x"78"),
  1209 => (x"c1",x"48",x"66",x"c4"),
  1210 => (x"58",x"a6",x"d0",x"88"),
  1211 => (x"c8",x"e3",x"87",x"c3"),
  1212 => (x"48",x"a6",x"d0",x"87"),
  1213 => (x"9c",x"74",x"78",x"c2"),
  1214 => (x"87",x"db",x"cd",x"02"),
  1215 => (x"c1",x"48",x"66",x"c8"),
  1216 => (x"03",x"a8",x"66",x"c8"),
  1217 => (x"dc",x"87",x"d0",x"cd"),
  1218 => (x"78",x"c0",x"48",x"a6"),
  1219 => (x"78",x"c0",x"80",x"e8"),
  1220 => (x"70",x"87",x"f6",x"e1"),
  1221 => (x"ac",x"d0",x"c1",x"4c"),
  1222 => (x"87",x"d7",x"c2",x"05"),
  1223 => (x"e4",x"7e",x"66",x"c4"),
  1224 => (x"49",x"70",x"87",x"da"),
  1225 => (x"e1",x"59",x"a6",x"c8"),
  1226 => (x"4c",x"70",x"87",x"df"),
  1227 => (x"05",x"ac",x"ec",x"c0"),
  1228 => (x"c8",x"87",x"eb",x"c1"),
  1229 => (x"91",x"cb",x"49",x"66"),
  1230 => (x"81",x"66",x"c0",x"c1"),
  1231 => (x"6a",x"4a",x"a1",x"c4"),
  1232 => (x"4a",x"a1",x"c8",x"4d"),
  1233 => (x"c1",x"52",x"66",x"c4"),
  1234 => (x"e0",x"79",x"cb",x"c4"),
  1235 => (x"4c",x"70",x"87",x"fb"),
  1236 => (x"87",x"d8",x"02",x"9c"),
  1237 => (x"02",x"ac",x"fb",x"c0"),
  1238 => (x"55",x"74",x"87",x"d2"),
  1239 => (x"70",x"87",x"ea",x"e0"),
  1240 => (x"c7",x"02",x"9c",x"4c"),
  1241 => (x"ac",x"fb",x"c0",x"87"),
  1242 => (x"87",x"ee",x"ff",x"05"),
  1243 => (x"c2",x"55",x"e0",x"c0"),
  1244 => (x"97",x"c0",x"55",x"c1"),
  1245 => (x"49",x"66",x"d8",x"7d"),
  1246 => (x"db",x"05",x"a9",x"6e"),
  1247 => (x"48",x"66",x"c8",x"87"),
  1248 => (x"04",x"a8",x"66",x"cc"),
  1249 => (x"66",x"c8",x"87",x"ca"),
  1250 => (x"cc",x"80",x"c1",x"48"),
  1251 => (x"87",x"c8",x"58",x"a6"),
  1252 => (x"c1",x"48",x"66",x"cc"),
  1253 => (x"58",x"a6",x"d0",x"88"),
  1254 => (x"87",x"ed",x"df",x"ff"),
  1255 => (x"d0",x"c1",x"4c",x"70"),
  1256 => (x"87",x"c8",x"05",x"ac"),
  1257 => (x"c1",x"48",x"66",x"d4"),
  1258 => (x"58",x"a6",x"d8",x"80"),
  1259 => (x"02",x"ac",x"d0",x"c1"),
  1260 => (x"c0",x"87",x"e9",x"fd"),
  1261 => (x"d8",x"48",x"a6",x"e0"),
  1262 => (x"66",x"c4",x"78",x"66"),
  1263 => (x"66",x"e0",x"c0",x"48"),
  1264 => (x"e4",x"c9",x"05",x"a8"),
  1265 => (x"a6",x"e4",x"c0",x"87"),
  1266 => (x"c4",x"78",x"c0",x"48"),
  1267 => (x"74",x"78",x"c0",x"80"),
  1268 => (x"88",x"fb",x"c0",x"48"),
  1269 => (x"02",x"6e",x"7e",x"70"),
  1270 => (x"6e",x"87",x"e7",x"c8"),
  1271 => (x"70",x"88",x"cb",x"48"),
  1272 => (x"c1",x"02",x"6e",x"7e"),
  1273 => (x"48",x"6e",x"87",x"cd"),
  1274 => (x"7e",x"70",x"88",x"c9"),
  1275 => (x"e9",x"c3",x"02",x"6e"),
  1276 => (x"c4",x"48",x"6e",x"87"),
  1277 => (x"6e",x"7e",x"70",x"88"),
  1278 => (x"6e",x"87",x"ce",x"02"),
  1279 => (x"70",x"88",x"c1",x"48"),
  1280 => (x"c3",x"02",x"6e",x"7e"),
  1281 => (x"f3",x"c7",x"87",x"d4"),
  1282 => (x"48",x"a6",x"dc",x"87"),
  1283 => (x"ff",x"78",x"f0",x"c0"),
  1284 => (x"70",x"87",x"f6",x"dd"),
  1285 => (x"ac",x"ec",x"c0",x"4c"),
  1286 => (x"87",x"c4",x"c0",x"02"),
  1287 => (x"5c",x"a6",x"e0",x"c0"),
  1288 => (x"02",x"ac",x"ec",x"c0"),
  1289 => (x"dd",x"ff",x"87",x"cd"),
  1290 => (x"4c",x"70",x"87",x"df"),
  1291 => (x"05",x"ac",x"ec",x"c0"),
  1292 => (x"c0",x"87",x"f3",x"ff"),
  1293 => (x"c0",x"02",x"ac",x"ec"),
  1294 => (x"dd",x"ff",x"87",x"c4"),
  1295 => (x"1e",x"c0",x"87",x"cb"),
  1296 => (x"66",x"d0",x"1e",x"ca"),
  1297 => (x"c1",x"91",x"cb",x"49"),
  1298 => (x"71",x"48",x"66",x"c8"),
  1299 => (x"58",x"a6",x"cc",x"80"),
  1300 => (x"c4",x"48",x"66",x"c8"),
  1301 => (x"58",x"a6",x"d0",x"80"),
  1302 => (x"49",x"bf",x"66",x"cc"),
  1303 => (x"87",x"ed",x"dd",x"ff"),
  1304 => (x"1e",x"de",x"1e",x"c1"),
  1305 => (x"49",x"bf",x"66",x"d4"),
  1306 => (x"87",x"e1",x"dd",x"ff"),
  1307 => (x"49",x"70",x"86",x"d0"),
  1308 => (x"c0",x"89",x"09",x"c0"),
  1309 => (x"c0",x"59",x"a6",x"ec"),
  1310 => (x"c0",x"48",x"66",x"e8"),
  1311 => (x"ee",x"c0",x"06",x"a8"),
  1312 => (x"66",x"e8",x"c0",x"87"),
  1313 => (x"03",x"a8",x"dd",x"48"),
  1314 => (x"c4",x"87",x"e4",x"c0"),
  1315 => (x"c0",x"49",x"bf",x"66"),
  1316 => (x"c0",x"81",x"66",x"e8"),
  1317 => (x"e8",x"c0",x"51",x"e0"),
  1318 => (x"81",x"c1",x"49",x"66"),
  1319 => (x"81",x"bf",x"66",x"c4"),
  1320 => (x"c0",x"51",x"c1",x"c2"),
  1321 => (x"c2",x"49",x"66",x"e8"),
  1322 => (x"bf",x"66",x"c4",x"81"),
  1323 => (x"6e",x"51",x"c0",x"81"),
  1324 => (x"ca",x"c3",x"c1",x"48"),
  1325 => (x"c8",x"49",x"6e",x"78"),
  1326 => (x"51",x"66",x"d0",x"81"),
  1327 => (x"81",x"c9",x"49",x"6e"),
  1328 => (x"6e",x"51",x"66",x"d4"),
  1329 => (x"dc",x"81",x"ca",x"49"),
  1330 => (x"66",x"d0",x"51",x"66"),
  1331 => (x"d4",x"80",x"c1",x"48"),
  1332 => (x"d8",x"48",x"58",x"a6"),
  1333 => (x"c4",x"78",x"c1",x"80"),
  1334 => (x"dd",x"ff",x"87",x"e8"),
  1335 => (x"49",x"70",x"87",x"de"),
  1336 => (x"59",x"a6",x"ec",x"c0"),
  1337 => (x"87",x"d4",x"dd",x"ff"),
  1338 => (x"e0",x"c0",x"49",x"70"),
  1339 => (x"66",x"dc",x"59",x"a6"),
  1340 => (x"a8",x"ec",x"c0",x"48"),
  1341 => (x"87",x"ca",x"c0",x"05"),
  1342 => (x"c0",x"48",x"a6",x"dc"),
  1343 => (x"c0",x"78",x"66",x"e8"),
  1344 => (x"da",x"ff",x"87",x"c4"),
  1345 => (x"66",x"c8",x"87",x"c3"),
  1346 => (x"c1",x"91",x"cb",x"49"),
  1347 => (x"71",x"48",x"66",x"c0"),
  1348 => (x"6e",x"7e",x"70",x"80"),
  1349 => (x"6e",x"82",x"c8",x"4a"),
  1350 => (x"c0",x"81",x"ca",x"49"),
  1351 => (x"dc",x"51",x"66",x"e8"),
  1352 => (x"81",x"c1",x"49",x"66"),
  1353 => (x"89",x"66",x"e8",x"c0"),
  1354 => (x"30",x"71",x"48",x"c1"),
  1355 => (x"89",x"c1",x"49",x"70"),
  1356 => (x"c2",x"7a",x"97",x"71"),
  1357 => (x"49",x"bf",x"f0",x"df"),
  1358 => (x"29",x"66",x"e8",x"c0"),
  1359 => (x"48",x"4a",x"6a",x"97"),
  1360 => (x"f0",x"c0",x"98",x"71"),
  1361 => (x"49",x"6e",x"58",x"a6"),
  1362 => (x"4d",x"69",x"81",x"c4"),
  1363 => (x"48",x"66",x"e0",x"c0"),
  1364 => (x"02",x"a8",x"66",x"c4"),
  1365 => (x"c4",x"87",x"c8",x"c0"),
  1366 => (x"78",x"c0",x"48",x"a6"),
  1367 => (x"c4",x"87",x"c5",x"c0"),
  1368 => (x"78",x"c1",x"48",x"a6"),
  1369 => (x"c0",x"1e",x"66",x"c4"),
  1370 => (x"49",x"75",x"1e",x"e0"),
  1371 => (x"87",x"dd",x"d9",x"ff"),
  1372 => (x"4c",x"70",x"86",x"c8"),
  1373 => (x"06",x"ac",x"b7",x"c0"),
  1374 => (x"74",x"87",x"d4",x"c1"),
  1375 => (x"49",x"e0",x"c0",x"85"),
  1376 => (x"4b",x"75",x"89",x"74"),
  1377 => (x"4a",x"d9",x"da",x"c1"),
  1378 => (x"db",x"ec",x"fe",x"71"),
  1379 => (x"c0",x"85",x"c2",x"87"),
  1380 => (x"c1",x"48",x"66",x"e4"),
  1381 => (x"a6",x"e8",x"c0",x"80"),
  1382 => (x"66",x"ec",x"c0",x"58"),
  1383 => (x"70",x"81",x"c1",x"49"),
  1384 => (x"c8",x"c0",x"02",x"a9"),
  1385 => (x"48",x"a6",x"c4",x"87"),
  1386 => (x"c5",x"c0",x"78",x"c0"),
  1387 => (x"48",x"a6",x"c4",x"87"),
  1388 => (x"66",x"c4",x"78",x"c1"),
  1389 => (x"49",x"a4",x"c2",x"1e"),
  1390 => (x"71",x"48",x"e0",x"c0"),
  1391 => (x"1e",x"49",x"70",x"88"),
  1392 => (x"d8",x"ff",x"49",x"75"),
  1393 => (x"86",x"c8",x"87",x"c7"),
  1394 => (x"01",x"a8",x"b7",x"c0"),
  1395 => (x"c0",x"87",x"c0",x"ff"),
  1396 => (x"c0",x"02",x"66",x"e4"),
  1397 => (x"49",x"6e",x"87",x"d1"),
  1398 => (x"e4",x"c0",x"81",x"c9"),
  1399 => (x"48",x"6e",x"51",x"66"),
  1400 => (x"78",x"db",x"c5",x"c1"),
  1401 => (x"6e",x"87",x"cc",x"c0"),
  1402 => (x"c2",x"81",x"c9",x"49"),
  1403 => (x"c1",x"48",x"6e",x"51"),
  1404 => (x"c0",x"78",x"cf",x"c6"),
  1405 => (x"c1",x"48",x"a6",x"e8"),
  1406 => (x"87",x"c6",x"c0",x"78"),
  1407 => (x"87",x"f9",x"d6",x"ff"),
  1408 => (x"e8",x"c0",x"4c",x"70"),
  1409 => (x"f5",x"c0",x"02",x"66"),
  1410 => (x"48",x"66",x"c8",x"87"),
  1411 => (x"04",x"a8",x"66",x"cc"),
  1412 => (x"c8",x"87",x"cb",x"c0"),
  1413 => (x"80",x"c1",x"48",x"66"),
  1414 => (x"c0",x"58",x"a6",x"cc"),
  1415 => (x"66",x"cc",x"87",x"e0"),
  1416 => (x"d0",x"88",x"c1",x"48"),
  1417 => (x"d5",x"c0",x"58",x"a6"),
  1418 => (x"ac",x"c6",x"c1",x"87"),
  1419 => (x"87",x"c8",x"c0",x"05"),
  1420 => (x"c1",x"48",x"66",x"d0"),
  1421 => (x"58",x"a6",x"d4",x"80"),
  1422 => (x"87",x"fd",x"d5",x"ff"),
  1423 => (x"66",x"d4",x"4c",x"70"),
  1424 => (x"d8",x"80",x"c1",x"48"),
  1425 => (x"9c",x"74",x"58",x"a6"),
  1426 => (x"87",x"cb",x"c0",x"02"),
  1427 => (x"c1",x"48",x"66",x"c8"),
  1428 => (x"04",x"a8",x"66",x"c8"),
  1429 => (x"ff",x"87",x"f0",x"f2"),
  1430 => (x"c8",x"87",x"d5",x"d5"),
  1431 => (x"a8",x"c7",x"48",x"66"),
  1432 => (x"87",x"e5",x"c0",x"03"),
  1433 => (x"48",x"c4",x"dc",x"c2"),
  1434 => (x"66",x"c8",x"78",x"c0"),
  1435 => (x"c1",x"91",x"cb",x"49"),
  1436 => (x"c4",x"81",x"66",x"c0"),
  1437 => (x"4a",x"6a",x"4a",x"a1"),
  1438 => (x"c8",x"79",x"52",x"c0"),
  1439 => (x"80",x"c1",x"48",x"66"),
  1440 => (x"c7",x"58",x"a6",x"cc"),
  1441 => (x"db",x"ff",x"04",x"a8"),
  1442 => (x"8e",x"d0",x"ff",x"87"),
  1443 => (x"87",x"e9",x"df",x"ff"),
  1444 => (x"64",x"61",x"6f",x"4c"),
  1445 => (x"20",x"2e",x"2a",x"20"),
  1446 => (x"00",x"20",x"3a",x"00"),
  1447 => (x"71",x"1e",x"73",x"1e"),
  1448 => (x"c6",x"02",x"9b",x"4b"),
  1449 => (x"c0",x"dc",x"c2",x"87"),
  1450 => (x"c7",x"78",x"c0",x"48"),
  1451 => (x"c0",x"dc",x"c2",x"1e"),
  1452 => (x"c1",x"1e",x"49",x"bf"),
  1453 => (x"c2",x"1e",x"c7",x"de"),
  1454 => (x"49",x"bf",x"e8",x"db"),
  1455 => (x"cc",x"87",x"f0",x"ed"),
  1456 => (x"e8",x"db",x"c2",x"86"),
  1457 => (x"ea",x"e9",x"49",x"bf"),
  1458 => (x"02",x"9b",x"73",x"87"),
  1459 => (x"de",x"c1",x"87",x"c8"),
  1460 => (x"e3",x"c0",x"49",x"c7"),
  1461 => (x"de",x"ff",x"87",x"fd"),
  1462 => (x"c1",x"1e",x"87",x"e3"),
  1463 => (x"c0",x"48",x"f3",x"dd"),
  1464 => (x"ea",x"df",x"c1",x"50"),
  1465 => (x"d9",x"ff",x"49",x"bf"),
  1466 => (x"48",x"c0",x"87",x"e1"),
  1467 => (x"c7",x"1e",x"4f",x"26"),
  1468 => (x"49",x"c1",x"87",x"df"),
  1469 => (x"fe",x"87",x"e5",x"fe"),
  1470 => (x"70",x"87",x"ee",x"ee"),
  1471 => (x"87",x"cd",x"02",x"98"),
  1472 => (x"87",x"c7",x"f6",x"fe"),
  1473 => (x"c4",x"02",x"98",x"70"),
  1474 => (x"c2",x"4a",x"c1",x"87"),
  1475 => (x"72",x"4a",x"c0",x"87"),
  1476 => (x"87",x"ce",x"05",x"9a"),
  1477 => (x"dc",x"c1",x"1e",x"c0"),
  1478 => (x"ef",x"c0",x"49",x"fe"),
  1479 => (x"86",x"c4",x"87",x"c3"),
  1480 => (x"1e",x"c0",x"87",x"fe"),
  1481 => (x"49",x"c9",x"dd",x"c1"),
  1482 => (x"87",x"f5",x"ee",x"c0"),
  1483 => (x"e9",x"fe",x"1e",x"c0"),
  1484 => (x"c0",x"49",x"70",x"87"),
  1485 => (x"c3",x"87",x"ea",x"ee"),
  1486 => (x"8e",x"f8",x"87",x"d6"),
  1487 => (x"44",x"53",x"4f",x"26"),
  1488 => (x"69",x"61",x"66",x"20"),
  1489 => (x"2e",x"64",x"65",x"6c"),
  1490 => (x"6f",x"6f",x"42",x"00"),
  1491 => (x"67",x"6e",x"69",x"74"),
  1492 => (x"00",x"2e",x"2e",x"2e"),
  1493 => (x"d6",x"e6",x"c0",x"1e"),
  1494 => (x"26",x"87",x"fa",x"87"),
  1495 => (x"dc",x"c2",x"1e",x"4f"),
  1496 => (x"78",x"c0",x"48",x"c0"),
  1497 => (x"48",x"e8",x"db",x"c2"),
  1498 => (x"c1",x"fe",x"78",x"c0"),
  1499 => (x"c0",x"87",x"e5",x"87"),
  1500 => (x"00",x"4f",x"26",x"48"),
  1501 => (x"00",x"00",x"01",x"00"),
  1502 => (x"45",x"20",x"80",x"00"),
  1503 => (x"00",x"74",x"69",x"78"),
  1504 => (x"61",x"42",x"20",x"80"),
  1505 => (x"0b",x"00",x"6b",x"63"),
  1506 => (x"14",x"00",x"00",x"11"),
  1507 => (x"00",x"00",x"00",x"27"),
  1508 => (x"11",x"0b",x"00",x"00"),
  1509 => (x"27",x"32",x"00",x"00"),
  1510 => (x"00",x"00",x"00",x"00"),
  1511 => (x"00",x"11",x"0b",x"00"),
  1512 => (x"00",x"27",x"50",x"00"),
  1513 => (x"00",x"00",x"00",x"00"),
  1514 => (x"00",x"00",x"11",x"0b"),
  1515 => (x"00",x"00",x"27",x"6e"),
  1516 => (x"0b",x"00",x"00",x"00"),
  1517 => (x"8c",x"00",x"00",x"11"),
  1518 => (x"00",x"00",x"00",x"27"),
  1519 => (x"11",x"0b",x"00",x"00"),
  1520 => (x"27",x"aa",x"00",x"00"),
  1521 => (x"00",x"00",x"00",x"00"),
  1522 => (x"00",x"11",x"0b",x"00"),
  1523 => (x"00",x"27",x"c8",x"00"),
  1524 => (x"00",x"00",x"00",x"00"),
  1525 => (x"00",x"00",x"11",x"0b"),
  1526 => (x"00",x"00",x"00",x"00"),
  1527 => (x"a0",x"00",x"00",x"00"),
  1528 => (x"00",x"00",x"00",x"11"),
  1529 => (x"00",x"00",x"00",x"00"),
  1530 => (x"17",x"ee",x"00",x"00"),
  1531 => (x"4f",x"42",x"00",x"00"),
  1532 => (x"20",x"20",x"54",x"4f"),
  1533 => (x"4f",x"52",x"20",x"20"),
  1534 => (x"fe",x"1e",x"00",x"4d"),
  1535 => (x"78",x"c0",x"48",x"f0"),
  1536 => (x"09",x"79",x"09",x"cd"),
  1537 => (x"1e",x"1e",x"4f",x"26"),
  1538 => (x"7e",x"bf",x"f0",x"fe"),
  1539 => (x"4f",x"26",x"26",x"48"),
  1540 => (x"48",x"f0",x"fe",x"1e"),
  1541 => (x"4f",x"26",x"78",x"c1"),
  1542 => (x"48",x"f0",x"fe",x"1e"),
  1543 => (x"4f",x"26",x"78",x"c0"),
  1544 => (x"c0",x"4a",x"71",x"1e"),
  1545 => (x"4f",x"26",x"52",x"52"),
  1546 => (x"5c",x"5b",x"5e",x"0e"),
  1547 => (x"86",x"f4",x"0e",x"5d"),
  1548 => (x"6d",x"97",x"4d",x"71"),
  1549 => (x"4c",x"a5",x"c1",x"7e"),
  1550 => (x"c8",x"48",x"6c",x"97"),
  1551 => (x"48",x"6e",x"58",x"a6"),
  1552 => (x"05",x"a8",x"66",x"c4"),
  1553 => (x"48",x"ff",x"87",x"c5"),
  1554 => (x"ff",x"87",x"e6",x"c0"),
  1555 => (x"a5",x"c2",x"87",x"ca"),
  1556 => (x"4b",x"6c",x"97",x"49"),
  1557 => (x"97",x"4b",x"a3",x"71"),
  1558 => (x"6c",x"97",x"4b",x"6b"),
  1559 => (x"c1",x"48",x"6e",x"7e"),
  1560 => (x"58",x"a6",x"c8",x"80"),
  1561 => (x"a6",x"cc",x"98",x"c7"),
  1562 => (x"7c",x"97",x"70",x"58"),
  1563 => (x"73",x"87",x"e1",x"fe"),
  1564 => (x"26",x"8e",x"f4",x"48"),
  1565 => (x"26",x"4c",x"26",x"4d"),
  1566 => (x"0e",x"4f",x"26",x"4b"),
  1567 => (x"0e",x"5c",x"5b",x"5e"),
  1568 => (x"4c",x"71",x"86",x"f4"),
  1569 => (x"c3",x"4a",x"66",x"d8"),
  1570 => (x"a4",x"c2",x"9a",x"ff"),
  1571 => (x"49",x"6c",x"97",x"4b"),
  1572 => (x"72",x"49",x"a1",x"73"),
  1573 => (x"7e",x"6c",x"97",x"51"),
  1574 => (x"80",x"c1",x"48",x"6e"),
  1575 => (x"c7",x"58",x"a6",x"c8"),
  1576 => (x"58",x"a6",x"cc",x"98"),
  1577 => (x"8e",x"f4",x"54",x"70"),
  1578 => (x"1e",x"87",x"ca",x"ff"),
  1579 => (x"87",x"e8",x"fd",x"1e"),
  1580 => (x"49",x"4a",x"bf",x"e0"),
  1581 => (x"99",x"c0",x"e0",x"c0"),
  1582 => (x"72",x"87",x"cb",x"02"),
  1583 => (x"e6",x"df",x"c2",x"1e"),
  1584 => (x"87",x"f7",x"fe",x"49"),
  1585 => (x"fd",x"fc",x"86",x"c4"),
  1586 => (x"fd",x"7e",x"70",x"87"),
  1587 => (x"26",x"26",x"87",x"c2"),
  1588 => (x"df",x"c2",x"1e",x"4f"),
  1589 => (x"c7",x"fd",x"49",x"e6"),
  1590 => (x"eb",x"e2",x"c1",x"87"),
  1591 => (x"87",x"da",x"fc",x"49"),
  1592 => (x"26",x"87",x"c7",x"c4"),
  1593 => (x"d0",x"ff",x"1e",x"4f"),
  1594 => (x"78",x"e1",x"c8",x"48"),
  1595 => (x"c5",x"48",x"d4",x"ff"),
  1596 => (x"02",x"66",x"c4",x"78"),
  1597 => (x"e0",x"c3",x"87",x"c3"),
  1598 => (x"02",x"66",x"c8",x"78"),
  1599 => (x"d4",x"ff",x"87",x"c6"),
  1600 => (x"78",x"f0",x"c3",x"48"),
  1601 => (x"71",x"48",x"d4",x"ff"),
  1602 => (x"48",x"d0",x"ff",x"78"),
  1603 => (x"c0",x"78",x"e1",x"c8"),
  1604 => (x"4f",x"26",x"78",x"e0"),
  1605 => (x"5c",x"5b",x"5e",x"0e"),
  1606 => (x"c2",x"4c",x"71",x"0e"),
  1607 => (x"fc",x"49",x"e6",x"df"),
  1608 => (x"4a",x"70",x"87",x"c6"),
  1609 => (x"04",x"aa",x"b7",x"c0"),
  1610 => (x"c3",x"87",x"e2",x"c2"),
  1611 => (x"c9",x"05",x"aa",x"f0"),
  1612 => (x"d9",x"e7",x"c1",x"87"),
  1613 => (x"c2",x"78",x"c1",x"48"),
  1614 => (x"e0",x"c3",x"87",x"c3"),
  1615 => (x"87",x"c9",x"05",x"aa"),
  1616 => (x"48",x"dd",x"e7",x"c1"),
  1617 => (x"f4",x"c1",x"78",x"c1"),
  1618 => (x"dd",x"e7",x"c1",x"87"),
  1619 => (x"87",x"c6",x"02",x"bf"),
  1620 => (x"4b",x"a2",x"c0",x"c2"),
  1621 => (x"4b",x"72",x"87",x"c2"),
  1622 => (x"d1",x"05",x"9c",x"74"),
  1623 => (x"d9",x"e7",x"c1",x"87"),
  1624 => (x"e7",x"c1",x"1e",x"bf"),
  1625 => (x"72",x"1e",x"bf",x"dd"),
  1626 => (x"87",x"f9",x"fd",x"49"),
  1627 => (x"e7",x"c1",x"86",x"c8"),
  1628 => (x"c0",x"02",x"bf",x"d9"),
  1629 => (x"49",x"73",x"87",x"e0"),
  1630 => (x"91",x"29",x"b7",x"c4"),
  1631 => (x"81",x"f9",x"e8",x"c1"),
  1632 => (x"9a",x"cf",x"4a",x"73"),
  1633 => (x"48",x"c1",x"92",x"c2"),
  1634 => (x"4a",x"70",x"30",x"72"),
  1635 => (x"48",x"72",x"ba",x"ff"),
  1636 => (x"79",x"70",x"98",x"69"),
  1637 => (x"49",x"73",x"87",x"db"),
  1638 => (x"91",x"29",x"b7",x"c4"),
  1639 => (x"81",x"f9",x"e8",x"c1"),
  1640 => (x"9a",x"cf",x"4a",x"73"),
  1641 => (x"48",x"c3",x"92",x"c2"),
  1642 => (x"4a",x"70",x"30",x"72"),
  1643 => (x"70",x"b0",x"69",x"48"),
  1644 => (x"dd",x"e7",x"c1",x"79"),
  1645 => (x"c1",x"78",x"c0",x"48"),
  1646 => (x"c0",x"48",x"d9",x"e7"),
  1647 => (x"e6",x"df",x"c2",x"78"),
  1648 => (x"87",x"e4",x"f9",x"49"),
  1649 => (x"b7",x"c0",x"4a",x"70"),
  1650 => (x"de",x"fd",x"03",x"aa"),
  1651 => (x"c2",x"48",x"c0",x"87"),
  1652 => (x"26",x"4d",x"26",x"87"),
  1653 => (x"26",x"4b",x"26",x"4c"),
  1654 => (x"00",x"00",x"00",x"4f"),
  1655 => (x"00",x"00",x"00",x"00"),
  1656 => (x"4a",x"71",x"1e",x"00"),
  1657 => (x"87",x"ec",x"fc",x"49"),
  1658 => (x"c0",x"1e",x"4f",x"26"),
  1659 => (x"c4",x"49",x"72",x"4a"),
  1660 => (x"f9",x"e8",x"c1",x"91"),
  1661 => (x"c1",x"79",x"c0",x"81"),
  1662 => (x"aa",x"b7",x"d0",x"82"),
  1663 => (x"26",x"87",x"ee",x"04"),
  1664 => (x"5b",x"5e",x"0e",x"4f"),
  1665 => (x"71",x"0e",x"5d",x"5c"),
  1666 => (x"87",x"cc",x"f8",x"4d"),
  1667 => (x"b7",x"c4",x"4a",x"75"),
  1668 => (x"e8",x"c1",x"92",x"2a"),
  1669 => (x"4c",x"75",x"82",x"f9"),
  1670 => (x"94",x"c2",x"9c",x"cf"),
  1671 => (x"74",x"4b",x"49",x"6a"),
  1672 => (x"c2",x"9b",x"c3",x"2b"),
  1673 => (x"70",x"30",x"74",x"48"),
  1674 => (x"74",x"bc",x"ff",x"4c"),
  1675 => (x"70",x"98",x"71",x"48"),
  1676 => (x"87",x"dc",x"f7",x"7a"),
  1677 => (x"d8",x"fe",x"48",x"73"),
  1678 => (x"00",x"00",x"00",x"87"),
  1679 => (x"00",x"00",x"00",x"00"),
  1680 => (x"00",x"00",x"00",x"00"),
  1681 => (x"00",x"00",x"00",x"00"),
  1682 => (x"00",x"00",x"00",x"00"),
  1683 => (x"00",x"00",x"00",x"00"),
  1684 => (x"00",x"00",x"00",x"00"),
  1685 => (x"00",x"00",x"00",x"00"),
  1686 => (x"00",x"00",x"00",x"00"),
  1687 => (x"00",x"00",x"00",x"00"),
  1688 => (x"00",x"00",x"00",x"00"),
  1689 => (x"00",x"00",x"00",x"00"),
  1690 => (x"00",x"00",x"00",x"00"),
  1691 => (x"00",x"00",x"00",x"00"),
  1692 => (x"00",x"00",x"00",x"00"),
  1693 => (x"00",x"00",x"00",x"00"),
  1694 => (x"d0",x"ff",x"1e",x"00"),
  1695 => (x"78",x"e1",x"c8",x"48"),
  1696 => (x"d4",x"ff",x"48",x"71"),
  1697 => (x"66",x"c4",x"78",x"08"),
  1698 => (x"08",x"d4",x"ff",x"48"),
  1699 => (x"1e",x"4f",x"26",x"78"),
  1700 => (x"66",x"c4",x"4a",x"71"),
  1701 => (x"49",x"72",x"1e",x"49"),
  1702 => (x"ff",x"87",x"de",x"ff"),
  1703 => (x"e0",x"c0",x"48",x"d0"),
  1704 => (x"4f",x"26",x"26",x"78"),
  1705 => (x"71",x"1e",x"73",x"1e"),
  1706 => (x"49",x"66",x"c8",x"4b"),
  1707 => (x"c1",x"4a",x"73",x"1e"),
  1708 => (x"ff",x"49",x"a2",x"e0"),
  1709 => (x"c4",x"26",x"87",x"d9"),
  1710 => (x"26",x"4d",x"26",x"87"),
  1711 => (x"26",x"4b",x"26",x"4c"),
  1712 => (x"d4",x"ff",x"1e",x"4f"),
  1713 => (x"7a",x"ff",x"c3",x"4a"),
  1714 => (x"c0",x"48",x"d0",x"ff"),
  1715 => (x"7a",x"de",x"78",x"e1"),
  1716 => (x"bf",x"f0",x"df",x"c2"),
  1717 => (x"c8",x"48",x"49",x"7a"),
  1718 => (x"71",x"7a",x"70",x"28"),
  1719 => (x"70",x"28",x"d0",x"48"),
  1720 => (x"d8",x"48",x"71",x"7a"),
  1721 => (x"ff",x"7a",x"70",x"28"),
  1722 => (x"e0",x"c0",x"48",x"d0"),
  1723 => (x"0e",x"4f",x"26",x"78"),
  1724 => (x"5d",x"5c",x"5b",x"5e"),
  1725 => (x"c2",x"4c",x"71",x"0e"),
  1726 => (x"4d",x"bf",x"f0",x"df"),
  1727 => (x"d0",x"2b",x"74",x"4b"),
  1728 => (x"83",x"c1",x"9b",x"66"),
  1729 => (x"04",x"ab",x"66",x"d4"),
  1730 => (x"4b",x"c0",x"87",x"c2"),
  1731 => (x"66",x"d0",x"4a",x"74"),
  1732 => (x"ff",x"31",x"72",x"49"),
  1733 => (x"73",x"99",x"75",x"b9"),
  1734 => (x"70",x"30",x"72",x"48"),
  1735 => (x"b0",x"71",x"48",x"4a"),
  1736 => (x"58",x"f4",x"df",x"c2"),
  1737 => (x"26",x"87",x"da",x"fe"),
  1738 => (x"26",x"4c",x"26",x"4d"),
  1739 => (x"1e",x"4f",x"26",x"4b"),
  1740 => (x"c8",x"48",x"d0",x"ff"),
  1741 => (x"48",x"71",x"78",x"c9"),
  1742 => (x"78",x"08",x"d4",x"ff"),
  1743 => (x"71",x"1e",x"4f",x"26"),
  1744 => (x"87",x"eb",x"49",x"4a"),
  1745 => (x"c8",x"48",x"d0",x"ff"),
  1746 => (x"1e",x"4f",x"26",x"78"),
  1747 => (x"4b",x"71",x"1e",x"73"),
  1748 => (x"bf",x"c0",x"e0",x"c2"),
  1749 => (x"c2",x"87",x"c3",x"02"),
  1750 => (x"d0",x"ff",x"87",x"eb"),
  1751 => (x"78",x"c9",x"c8",x"48"),
  1752 => (x"e0",x"c0",x"49",x"73"),
  1753 => (x"48",x"d4",x"ff",x"b1"),
  1754 => (x"df",x"c2",x"78",x"71"),
  1755 => (x"78",x"c0",x"48",x"f4"),
  1756 => (x"c5",x"02",x"66",x"c8"),
  1757 => (x"49",x"ff",x"c3",x"87"),
  1758 => (x"49",x"c0",x"87",x"c2"),
  1759 => (x"59",x"fc",x"df",x"c2"),
  1760 => (x"c6",x"02",x"66",x"cc"),
  1761 => (x"d5",x"d5",x"c5",x"87"),
  1762 => (x"cf",x"87",x"c4",x"4a"),
  1763 => (x"c2",x"4a",x"ff",x"ff"),
  1764 => (x"c2",x"5a",x"c0",x"e0"),
  1765 => (x"c1",x"48",x"c0",x"e0"),
  1766 => (x"26",x"87",x"c4",x"78"),
  1767 => (x"26",x"4c",x"26",x"4d"),
  1768 => (x"0e",x"4f",x"26",x"4b"),
  1769 => (x"5d",x"5c",x"5b",x"5e"),
  1770 => (x"c2",x"4a",x"71",x"0e"),
  1771 => (x"4c",x"bf",x"fc",x"df"),
  1772 => (x"cb",x"02",x"9a",x"72"),
  1773 => (x"91",x"c8",x"49",x"87"),
  1774 => (x"4b",x"c1",x"ed",x"c1"),
  1775 => (x"87",x"c4",x"83",x"71"),
  1776 => (x"4b",x"c1",x"f1",x"c1"),
  1777 => (x"49",x"13",x"4d",x"c0"),
  1778 => (x"df",x"c2",x"99",x"74"),
  1779 => (x"ff",x"b9",x"bf",x"f8"),
  1780 => (x"78",x"71",x"48",x"d4"),
  1781 => (x"85",x"2c",x"b7",x"c1"),
  1782 => (x"04",x"ad",x"b7",x"c8"),
  1783 => (x"df",x"c2",x"87",x"e8"),
  1784 => (x"c8",x"48",x"bf",x"f4"),
  1785 => (x"f8",x"df",x"c2",x"80"),
  1786 => (x"87",x"ef",x"fe",x"58"),
  1787 => (x"71",x"1e",x"73",x"1e"),
  1788 => (x"9a",x"4a",x"13",x"4b"),
  1789 => (x"72",x"87",x"cb",x"02"),
  1790 => (x"87",x"e7",x"fe",x"49"),
  1791 => (x"05",x"9a",x"4a",x"13"),
  1792 => (x"da",x"fe",x"87",x"f5"),
  1793 => (x"df",x"c2",x"1e",x"87"),
  1794 => (x"c2",x"49",x"bf",x"f4"),
  1795 => (x"c1",x"48",x"f4",x"df"),
  1796 => (x"c0",x"c4",x"78",x"a1"),
  1797 => (x"db",x"03",x"a9",x"b7"),
  1798 => (x"48",x"d4",x"ff",x"87"),
  1799 => (x"bf",x"f8",x"df",x"c2"),
  1800 => (x"f4",x"df",x"c2",x"78"),
  1801 => (x"df",x"c2",x"49",x"bf"),
  1802 => (x"a1",x"c1",x"48",x"f4"),
  1803 => (x"b7",x"c0",x"c4",x"78"),
  1804 => (x"87",x"e5",x"04",x"a9"),
  1805 => (x"c8",x"48",x"d0",x"ff"),
  1806 => (x"c0",x"e0",x"c2",x"78"),
  1807 => (x"26",x"78",x"c0",x"48"),
  1808 => (x"00",x"00",x"00",x"4f"),
  1809 => (x"00",x"00",x"00",x"00"),
  1810 => (x"00",x"00",x"00",x"00"),
  1811 => (x"00",x"00",x"5f",x"5f"),
  1812 => (x"03",x"03",x"00",x"00"),
  1813 => (x"00",x"03",x"03",x"00"),
  1814 => (x"7f",x"7f",x"14",x"00"),
  1815 => (x"14",x"7f",x"7f",x"14"),
  1816 => (x"2e",x"24",x"00",x"00"),
  1817 => (x"12",x"3a",x"6b",x"6b"),
  1818 => (x"36",x"6a",x"4c",x"00"),
  1819 => (x"32",x"56",x"6c",x"18"),
  1820 => (x"4f",x"7e",x"30",x"00"),
  1821 => (x"68",x"3a",x"77",x"59"),
  1822 => (x"04",x"00",x"00",x"40"),
  1823 => (x"00",x"00",x"03",x"07"),
  1824 => (x"1c",x"00",x"00",x"00"),
  1825 => (x"00",x"41",x"63",x"3e"),
  1826 => (x"41",x"00",x"00",x"00"),
  1827 => (x"00",x"1c",x"3e",x"63"),
  1828 => (x"3e",x"2a",x"08",x"00"),
  1829 => (x"2a",x"3e",x"1c",x"1c"),
  1830 => (x"08",x"08",x"00",x"08"),
  1831 => (x"08",x"08",x"3e",x"3e"),
  1832 => (x"80",x"00",x"00",x"00"),
  1833 => (x"00",x"00",x"60",x"e0"),
  1834 => (x"08",x"08",x"00",x"00"),
  1835 => (x"08",x"08",x"08",x"08"),
  1836 => (x"00",x"00",x"00",x"00"),
  1837 => (x"00",x"00",x"60",x"60"),
  1838 => (x"30",x"60",x"40",x"00"),
  1839 => (x"03",x"06",x"0c",x"18"),
  1840 => (x"7f",x"3e",x"00",x"01"),
  1841 => (x"3e",x"7f",x"4d",x"59"),
  1842 => (x"06",x"04",x"00",x"00"),
  1843 => (x"00",x"00",x"7f",x"7f"),
  1844 => (x"63",x"42",x"00",x"00"),
  1845 => (x"46",x"4f",x"59",x"71"),
  1846 => (x"63",x"22",x"00",x"00"),
  1847 => (x"36",x"7f",x"49",x"49"),
  1848 => (x"16",x"1c",x"18",x"00"),
  1849 => (x"10",x"7f",x"7f",x"13"),
  1850 => (x"67",x"27",x"00",x"00"),
  1851 => (x"39",x"7d",x"45",x"45"),
  1852 => (x"7e",x"3c",x"00",x"00"),
  1853 => (x"30",x"79",x"49",x"4b"),
  1854 => (x"01",x"01",x"00",x"00"),
  1855 => (x"07",x"0f",x"79",x"71"),
  1856 => (x"7f",x"36",x"00",x"00"),
  1857 => (x"36",x"7f",x"49",x"49"),
  1858 => (x"4f",x"06",x"00",x"00"),
  1859 => (x"1e",x"3f",x"69",x"49"),
  1860 => (x"00",x"00",x"00",x"00"),
  1861 => (x"00",x"00",x"66",x"66"),
  1862 => (x"80",x"00",x"00",x"00"),
  1863 => (x"00",x"00",x"66",x"e6"),
  1864 => (x"08",x"08",x"00",x"00"),
  1865 => (x"22",x"22",x"14",x"14"),
  1866 => (x"14",x"14",x"00",x"00"),
  1867 => (x"14",x"14",x"14",x"14"),
  1868 => (x"22",x"22",x"00",x"00"),
  1869 => (x"08",x"08",x"14",x"14"),
  1870 => (x"03",x"02",x"00",x"00"),
  1871 => (x"06",x"0f",x"59",x"51"),
  1872 => (x"41",x"7f",x"3e",x"00"),
  1873 => (x"1e",x"1f",x"55",x"5d"),
  1874 => (x"7f",x"7e",x"00",x"00"),
  1875 => (x"7e",x"7f",x"09",x"09"),
  1876 => (x"7f",x"7f",x"00",x"00"),
  1877 => (x"36",x"7f",x"49",x"49"),
  1878 => (x"3e",x"1c",x"00",x"00"),
  1879 => (x"41",x"41",x"41",x"63"),
  1880 => (x"7f",x"7f",x"00",x"00"),
  1881 => (x"1c",x"3e",x"63",x"41"),
  1882 => (x"7f",x"7f",x"00",x"00"),
  1883 => (x"41",x"41",x"49",x"49"),
  1884 => (x"7f",x"7f",x"00",x"00"),
  1885 => (x"01",x"01",x"09",x"09"),
  1886 => (x"7f",x"3e",x"00",x"00"),
  1887 => (x"7a",x"7b",x"49",x"41"),
  1888 => (x"7f",x"7f",x"00",x"00"),
  1889 => (x"7f",x"7f",x"08",x"08"),
  1890 => (x"41",x"00",x"00",x"00"),
  1891 => (x"00",x"41",x"7f",x"7f"),
  1892 => (x"60",x"20",x"00",x"00"),
  1893 => (x"3f",x"7f",x"40",x"40"),
  1894 => (x"08",x"7f",x"7f",x"00"),
  1895 => (x"41",x"63",x"36",x"1c"),
  1896 => (x"7f",x"7f",x"00",x"00"),
  1897 => (x"40",x"40",x"40",x"40"),
  1898 => (x"06",x"7f",x"7f",x"00"),
  1899 => (x"7f",x"7f",x"06",x"0c"),
  1900 => (x"06",x"7f",x"7f",x"00"),
  1901 => (x"7f",x"7f",x"18",x"0c"),
  1902 => (x"7f",x"3e",x"00",x"00"),
  1903 => (x"3e",x"7f",x"41",x"41"),
  1904 => (x"7f",x"7f",x"00",x"00"),
  1905 => (x"06",x"0f",x"09",x"09"),
  1906 => (x"41",x"7f",x"3e",x"00"),
  1907 => (x"40",x"7e",x"7f",x"61"),
  1908 => (x"7f",x"7f",x"00",x"00"),
  1909 => (x"66",x"7f",x"19",x"09"),
  1910 => (x"6f",x"26",x"00",x"00"),
  1911 => (x"32",x"7b",x"59",x"4d"),
  1912 => (x"01",x"01",x"00",x"00"),
  1913 => (x"01",x"01",x"7f",x"7f"),
  1914 => (x"7f",x"3f",x"00",x"00"),
  1915 => (x"3f",x"7f",x"40",x"40"),
  1916 => (x"3f",x"0f",x"00",x"00"),
  1917 => (x"0f",x"3f",x"70",x"70"),
  1918 => (x"30",x"7f",x"7f",x"00"),
  1919 => (x"7f",x"7f",x"30",x"18"),
  1920 => (x"36",x"63",x"41",x"00"),
  1921 => (x"63",x"36",x"1c",x"1c"),
  1922 => (x"06",x"03",x"01",x"41"),
  1923 => (x"03",x"06",x"7c",x"7c"),
  1924 => (x"59",x"71",x"61",x"01"),
  1925 => (x"41",x"43",x"47",x"4d"),
  1926 => (x"7f",x"00",x"00",x"00"),
  1927 => (x"00",x"41",x"41",x"7f"),
  1928 => (x"06",x"03",x"01",x"00"),
  1929 => (x"60",x"30",x"18",x"0c"),
  1930 => (x"41",x"00",x"00",x"40"),
  1931 => (x"00",x"7f",x"7f",x"41"),
  1932 => (x"06",x"0c",x"08",x"00"),
  1933 => (x"08",x"0c",x"06",x"03"),
  1934 => (x"80",x"80",x"80",x"00"),
  1935 => (x"80",x"80",x"80",x"80"),
  1936 => (x"00",x"00",x"00",x"00"),
  1937 => (x"00",x"04",x"07",x"03"),
  1938 => (x"74",x"20",x"00",x"00"),
  1939 => (x"78",x"7c",x"54",x"54"),
  1940 => (x"7f",x"7f",x"00",x"00"),
  1941 => (x"38",x"7c",x"44",x"44"),
  1942 => (x"7c",x"38",x"00",x"00"),
  1943 => (x"00",x"44",x"44",x"44"),
  1944 => (x"7c",x"38",x"00",x"00"),
  1945 => (x"7f",x"7f",x"44",x"44"),
  1946 => (x"7c",x"38",x"00",x"00"),
  1947 => (x"18",x"5c",x"54",x"54"),
  1948 => (x"7e",x"04",x"00",x"00"),
  1949 => (x"00",x"05",x"05",x"7f"),
  1950 => (x"bc",x"18",x"00",x"00"),
  1951 => (x"7c",x"fc",x"a4",x"a4"),
  1952 => (x"7f",x"7f",x"00",x"00"),
  1953 => (x"78",x"7c",x"04",x"04"),
  1954 => (x"00",x"00",x"00",x"00"),
  1955 => (x"00",x"40",x"7d",x"3d"),
  1956 => (x"80",x"80",x"00",x"00"),
  1957 => (x"00",x"7d",x"fd",x"80"),
  1958 => (x"7f",x"7f",x"00",x"00"),
  1959 => (x"44",x"6c",x"38",x"10"),
  1960 => (x"00",x"00",x"00",x"00"),
  1961 => (x"00",x"40",x"7f",x"3f"),
  1962 => (x"0c",x"7c",x"7c",x"00"),
  1963 => (x"78",x"7c",x"0c",x"18"),
  1964 => (x"7c",x"7c",x"00",x"00"),
  1965 => (x"78",x"7c",x"04",x"04"),
  1966 => (x"7c",x"38",x"00",x"00"),
  1967 => (x"38",x"7c",x"44",x"44"),
  1968 => (x"fc",x"fc",x"00",x"00"),
  1969 => (x"18",x"3c",x"24",x"24"),
  1970 => (x"3c",x"18",x"00",x"00"),
  1971 => (x"fc",x"fc",x"24",x"24"),
  1972 => (x"7c",x"7c",x"00",x"00"),
  1973 => (x"08",x"0c",x"04",x"04"),
  1974 => (x"5c",x"48",x"00",x"00"),
  1975 => (x"20",x"74",x"54",x"54"),
  1976 => (x"3f",x"04",x"00",x"00"),
  1977 => (x"00",x"44",x"44",x"7f"),
  1978 => (x"7c",x"3c",x"00",x"00"),
  1979 => (x"7c",x"7c",x"40",x"40"),
  1980 => (x"3c",x"1c",x"00",x"00"),
  1981 => (x"1c",x"3c",x"60",x"60"),
  1982 => (x"60",x"7c",x"3c",x"00"),
  1983 => (x"3c",x"7c",x"60",x"30"),
  1984 => (x"38",x"6c",x"44",x"00"),
  1985 => (x"44",x"6c",x"38",x"10"),
  1986 => (x"bc",x"1c",x"00",x"00"),
  1987 => (x"1c",x"3c",x"60",x"e0"),
  1988 => (x"64",x"44",x"00",x"00"),
  1989 => (x"44",x"4c",x"5c",x"74"),
  1990 => (x"08",x"08",x"00",x"00"),
  1991 => (x"41",x"41",x"77",x"3e"),
  1992 => (x"00",x"00",x"00",x"00"),
  1993 => (x"00",x"00",x"7f",x"7f"),
  1994 => (x"41",x"41",x"00",x"00"),
  1995 => (x"08",x"08",x"3e",x"77"),
  1996 => (x"01",x"01",x"02",x"00"),
  1997 => (x"01",x"02",x"02",x"03"),
  1998 => (x"7f",x"7f",x"7f",x"00"),
  1999 => (x"7f",x"7f",x"7f",x"7f"),
  2000 => (x"1c",x"08",x"08",x"00"),
  2001 => (x"7f",x"3e",x"3e",x"1c"),
  2002 => (x"3e",x"7f",x"7f",x"7f"),
  2003 => (x"08",x"1c",x"1c",x"3e"),
  2004 => (x"18",x"10",x"00",x"08"),
  2005 => (x"10",x"18",x"7c",x"7c"),
  2006 => (x"30",x"10",x"00",x"00"),
  2007 => (x"10",x"30",x"7c",x"7c"),
  2008 => (x"60",x"30",x"10",x"00"),
  2009 => (x"06",x"1e",x"78",x"60"),
  2010 => (x"3c",x"66",x"42",x"00"),
  2011 => (x"42",x"66",x"3c",x"18"),
  2012 => (x"6a",x"38",x"78",x"00"),
  2013 => (x"38",x"6c",x"c6",x"c2"),
  2014 => (x"00",x"00",x"60",x"00"),
  2015 => (x"60",x"00",x"00",x"60"),
  2016 => (x"5b",x"5e",x"0e",x"00"),
  2017 => (x"1e",x"0e",x"5d",x"5c"),
  2018 => (x"e0",x"c2",x"4c",x"71"),
  2019 => (x"c0",x"4d",x"bf",x"d1"),
  2020 => (x"74",x"1e",x"c0",x"4b"),
  2021 => (x"87",x"c7",x"02",x"ab"),
  2022 => (x"c0",x"48",x"a6",x"c4"),
  2023 => (x"c4",x"87",x"c5",x"78"),
  2024 => (x"78",x"c1",x"48",x"a6"),
  2025 => (x"73",x"1e",x"66",x"c4"),
  2026 => (x"87",x"df",x"ee",x"49"),
  2027 => (x"e0",x"c0",x"86",x"c8"),
  2028 => (x"87",x"ef",x"ef",x"49"),
  2029 => (x"6a",x"4a",x"a5",x"c4"),
  2030 => (x"87",x"f0",x"f0",x"49"),
  2031 => (x"cb",x"87",x"c6",x"f1"),
  2032 => (x"c8",x"83",x"c1",x"85"),
  2033 => (x"ff",x"04",x"ab",x"b7"),
  2034 => (x"26",x"26",x"87",x"c7"),
  2035 => (x"26",x"4c",x"26",x"4d"),
  2036 => (x"1e",x"4f",x"26",x"4b"),
  2037 => (x"e0",x"c2",x"4a",x"71"),
  2038 => (x"e0",x"c2",x"5a",x"d5"),
  2039 => (x"78",x"c7",x"48",x"d5"),
  2040 => (x"87",x"dd",x"fe",x"49"),
  2041 => (x"73",x"1e",x"4f",x"26"),
  2042 => (x"c0",x"4a",x"71",x"1e"),
  2043 => (x"d3",x"03",x"aa",x"b7"),
  2044 => (x"f6",x"cc",x"c2",x"87"),
  2045 => (x"87",x"c4",x"05",x"bf"),
  2046 => (x"87",x"c2",x"4b",x"c1"),
  2047 => (x"cc",x"c2",x"4b",x"c0"),
  2048 => (x"87",x"c4",x"5b",x"fa"),
  2049 => (x"5a",x"fa",x"cc",x"c2"),
  2050 => (x"bf",x"f6",x"cc",x"c2"),
  2051 => (x"c1",x"9a",x"c1",x"4a"),
  2052 => (x"ec",x"49",x"a2",x"c0"),
  2053 => (x"48",x"fc",x"87",x"e8"),
  2054 => (x"bf",x"f6",x"cc",x"c2"),
  2055 => (x"87",x"ef",x"fe",x"78"),
  2056 => (x"c4",x"4a",x"71",x"1e"),
  2057 => (x"49",x"72",x"1e",x"66"),
  2058 => (x"26",x"87",x"f9",x"e9"),
  2059 => (x"c2",x"1e",x"4f",x"26"),
  2060 => (x"49",x"bf",x"f6",x"cc"),
  2061 => (x"c2",x"87",x"ea",x"e6"),
  2062 => (x"e8",x"48",x"c9",x"e0"),
  2063 => (x"e0",x"c2",x"78",x"bf"),
  2064 => (x"bf",x"ec",x"48",x"c5"),
  2065 => (x"c9",x"e0",x"c2",x"78"),
  2066 => (x"c3",x"49",x"4a",x"bf"),
  2067 => (x"b7",x"c8",x"99",x"ff"),
  2068 => (x"71",x"48",x"72",x"2a"),
  2069 => (x"d1",x"e0",x"c2",x"b0"),
  2070 => (x"0e",x"4f",x"26",x"58"),
  2071 => (x"5d",x"5c",x"5b",x"5e"),
  2072 => (x"ff",x"4b",x"71",x"0e"),
  2073 => (x"e0",x"c2",x"87",x"c8"),
  2074 => (x"50",x"c0",x"48",x"c4"),
  2075 => (x"d0",x"e6",x"49",x"73"),
  2076 => (x"4c",x"49",x"70",x"87"),
  2077 => (x"ee",x"cb",x"9c",x"c2"),
  2078 => (x"87",x"c2",x"cb",x"49"),
  2079 => (x"c2",x"4d",x"49",x"70"),
  2080 => (x"bf",x"97",x"c4",x"e0"),
  2081 => (x"87",x"e2",x"c1",x"05"),
  2082 => (x"c2",x"49",x"66",x"d0"),
  2083 => (x"99",x"bf",x"cd",x"e0"),
  2084 => (x"d4",x"87",x"d6",x"05"),
  2085 => (x"e0",x"c2",x"49",x"66"),
  2086 => (x"05",x"99",x"bf",x"c5"),
  2087 => (x"49",x"73",x"87",x"cb"),
  2088 => (x"70",x"87",x"de",x"e5"),
  2089 => (x"c1",x"c1",x"02",x"98"),
  2090 => (x"fe",x"4c",x"c1",x"87"),
  2091 => (x"49",x"75",x"87",x"c0"),
  2092 => (x"70",x"87",x"d7",x"ca"),
  2093 => (x"87",x"c6",x"02",x"98"),
  2094 => (x"48",x"c4",x"e0",x"c2"),
  2095 => (x"e0",x"c2",x"50",x"c1"),
  2096 => (x"05",x"bf",x"97",x"c4"),
  2097 => (x"c2",x"87",x"e3",x"c0"),
  2098 => (x"49",x"bf",x"cd",x"e0"),
  2099 => (x"05",x"99",x"66",x"d0"),
  2100 => (x"c2",x"87",x"d6",x"ff"),
  2101 => (x"49",x"bf",x"c5",x"e0"),
  2102 => (x"05",x"99",x"66",x"d4"),
  2103 => (x"73",x"87",x"ca",x"ff"),
  2104 => (x"87",x"dd",x"e4",x"49"),
  2105 => (x"fe",x"05",x"98",x"70"),
  2106 => (x"48",x"74",x"87",x"ff"),
  2107 => (x"0e",x"87",x"dc",x"fb"),
  2108 => (x"5d",x"5c",x"5b",x"5e"),
  2109 => (x"c0",x"86",x"f4",x"0e"),
  2110 => (x"bf",x"ec",x"4c",x"4d"),
  2111 => (x"48",x"a6",x"c4",x"7e"),
  2112 => (x"bf",x"d1",x"e0",x"c2"),
  2113 => (x"c0",x"1e",x"c1",x"78"),
  2114 => (x"fd",x"49",x"c7",x"1e"),
  2115 => (x"86",x"c8",x"87",x"cd"),
  2116 => (x"cd",x"02",x"98",x"70"),
  2117 => (x"fb",x"49",x"ff",x"87"),
  2118 => (x"da",x"c1",x"87",x"cc"),
  2119 => (x"87",x"e1",x"e3",x"49"),
  2120 => (x"e0",x"c2",x"4d",x"c1"),
  2121 => (x"02",x"bf",x"97",x"c4"),
  2122 => (x"f6",x"c8",x"87",x"c3"),
  2123 => (x"c9",x"e0",x"c2",x"87"),
  2124 => (x"cc",x"c2",x"4b",x"bf"),
  2125 => (x"c0",x"05",x"bf",x"f6"),
  2126 => (x"fd",x"c3",x"87",x"e9"),
  2127 => (x"87",x"c1",x"e3",x"49"),
  2128 => (x"e2",x"49",x"fa",x"c3"),
  2129 => (x"49",x"73",x"87",x"fb"),
  2130 => (x"71",x"99",x"ff",x"c3"),
  2131 => (x"fb",x"49",x"c0",x"1e"),
  2132 => (x"49",x"73",x"87",x"ce"),
  2133 => (x"71",x"29",x"b7",x"c8"),
  2134 => (x"fb",x"49",x"c1",x"1e"),
  2135 => (x"86",x"c8",x"87",x"c2"),
  2136 => (x"c2",x"87",x"f9",x"c5"),
  2137 => (x"4b",x"bf",x"cd",x"e0"),
  2138 => (x"87",x"dd",x"02",x"9b"),
  2139 => (x"bf",x"f2",x"cc",x"c2"),
  2140 => (x"87",x"d6",x"c7",x"49"),
  2141 => (x"c4",x"05",x"98",x"70"),
  2142 => (x"d2",x"4b",x"c0",x"87"),
  2143 => (x"49",x"e0",x"c2",x"87"),
  2144 => (x"c2",x"87",x"fb",x"c6"),
  2145 => (x"c6",x"58",x"f6",x"cc"),
  2146 => (x"f2",x"cc",x"c2",x"87"),
  2147 => (x"73",x"78",x"c0",x"48"),
  2148 => (x"05",x"99",x"c2",x"49"),
  2149 => (x"eb",x"c3",x"87",x"cd"),
  2150 => (x"87",x"e5",x"e1",x"49"),
  2151 => (x"99",x"c2",x"49",x"70"),
  2152 => (x"fb",x"87",x"c2",x"02"),
  2153 => (x"c1",x"49",x"73",x"4c"),
  2154 => (x"87",x"cd",x"05",x"99"),
  2155 => (x"e1",x"49",x"f4",x"c3"),
  2156 => (x"49",x"70",x"87",x"cf"),
  2157 => (x"c2",x"02",x"99",x"c2"),
  2158 => (x"73",x"4c",x"fa",x"87"),
  2159 => (x"05",x"99",x"c8",x"49"),
  2160 => (x"f5",x"c3",x"87",x"cd"),
  2161 => (x"87",x"f9",x"e0",x"49"),
  2162 => (x"99",x"c2",x"49",x"70"),
  2163 => (x"c2",x"87",x"d4",x"02"),
  2164 => (x"02",x"bf",x"d5",x"e0"),
  2165 => (x"c1",x"48",x"87",x"c9"),
  2166 => (x"d9",x"e0",x"c2",x"88"),
  2167 => (x"ff",x"87",x"c2",x"58"),
  2168 => (x"73",x"4d",x"c1",x"4c"),
  2169 => (x"05",x"99",x"c4",x"49"),
  2170 => (x"f2",x"c3",x"87",x"cd"),
  2171 => (x"87",x"d1",x"e0",x"49"),
  2172 => (x"99",x"c2",x"49",x"70"),
  2173 => (x"c2",x"87",x"db",x"02"),
  2174 => (x"7e",x"bf",x"d5",x"e0"),
  2175 => (x"a8",x"b7",x"c7",x"48"),
  2176 => (x"6e",x"87",x"cb",x"03"),
  2177 => (x"c2",x"80",x"c1",x"48"),
  2178 => (x"c0",x"58",x"d9",x"e0"),
  2179 => (x"4c",x"fe",x"87",x"c2"),
  2180 => (x"fd",x"c3",x"4d",x"c1"),
  2181 => (x"e8",x"df",x"ff",x"49"),
  2182 => (x"c2",x"49",x"70",x"87"),
  2183 => (x"87",x"d5",x"02",x"99"),
  2184 => (x"bf",x"d5",x"e0",x"c2"),
  2185 => (x"87",x"c9",x"c0",x"02"),
  2186 => (x"48",x"d5",x"e0",x"c2"),
  2187 => (x"c2",x"c0",x"78",x"c0"),
  2188 => (x"c1",x"4c",x"fd",x"87"),
  2189 => (x"49",x"fa",x"c3",x"4d"),
  2190 => (x"87",x"c5",x"df",x"ff"),
  2191 => (x"99",x"c2",x"49",x"70"),
  2192 => (x"c2",x"87",x"d9",x"02"),
  2193 => (x"48",x"bf",x"d5",x"e0"),
  2194 => (x"03",x"a8",x"b7",x"c7"),
  2195 => (x"c2",x"87",x"c9",x"c0"),
  2196 => (x"c7",x"48",x"d5",x"e0"),
  2197 => (x"87",x"c2",x"c0",x"78"),
  2198 => (x"4d",x"c1",x"4c",x"fc"),
  2199 => (x"03",x"ac",x"b7",x"c0"),
  2200 => (x"c4",x"87",x"d1",x"c0"),
  2201 => (x"d8",x"c1",x"4a",x"66"),
  2202 => (x"c0",x"02",x"6a",x"82"),
  2203 => (x"4b",x"6a",x"87",x"c6"),
  2204 => (x"0f",x"73",x"49",x"74"),
  2205 => (x"f0",x"c3",x"1e",x"c0"),
  2206 => (x"49",x"da",x"c1",x"1e"),
  2207 => (x"c8",x"87",x"dc",x"f7"),
  2208 => (x"02",x"98",x"70",x"86"),
  2209 => (x"c8",x"87",x"e2",x"c0"),
  2210 => (x"e0",x"c2",x"48",x"a6"),
  2211 => (x"c8",x"78",x"bf",x"d5"),
  2212 => (x"91",x"cb",x"49",x"66"),
  2213 => (x"71",x"48",x"66",x"c4"),
  2214 => (x"6e",x"7e",x"70",x"80"),
  2215 => (x"c8",x"c0",x"02",x"bf"),
  2216 => (x"4b",x"bf",x"6e",x"87"),
  2217 => (x"73",x"49",x"66",x"c8"),
  2218 => (x"02",x"9d",x"75",x"0f"),
  2219 => (x"c2",x"87",x"c8",x"c0"),
  2220 => (x"49",x"bf",x"d5",x"e0"),
  2221 => (x"c2",x"87",x"ca",x"f3"),
  2222 => (x"02",x"bf",x"fa",x"cc"),
  2223 => (x"49",x"87",x"dd",x"c0"),
  2224 => (x"70",x"87",x"c7",x"c2"),
  2225 => (x"d3",x"c0",x"02",x"98"),
  2226 => (x"d5",x"e0",x"c2",x"87"),
  2227 => (x"f0",x"f2",x"49",x"bf"),
  2228 => (x"f4",x"49",x"c0",x"87"),
  2229 => (x"cc",x"c2",x"87",x"d0"),
  2230 => (x"78",x"c0",x"48",x"fa"),
  2231 => (x"ea",x"f3",x"8e",x"f4"),
  2232 => (x"5b",x"5e",x"0e",x"87"),
  2233 => (x"1e",x"0e",x"5d",x"5c"),
  2234 => (x"e0",x"c2",x"4c",x"71"),
  2235 => (x"c1",x"49",x"bf",x"d1"),
  2236 => (x"c1",x"4d",x"a1",x"cd"),
  2237 => (x"7e",x"69",x"81",x"d1"),
  2238 => (x"cf",x"02",x"9c",x"74"),
  2239 => (x"4b",x"a5",x"c4",x"87"),
  2240 => (x"e0",x"c2",x"7b",x"74"),
  2241 => (x"f3",x"49",x"bf",x"d1"),
  2242 => (x"7b",x"6e",x"87",x"c9"),
  2243 => (x"c4",x"05",x"9c",x"74"),
  2244 => (x"c2",x"4b",x"c0",x"87"),
  2245 => (x"73",x"4b",x"c1",x"87"),
  2246 => (x"87",x"ca",x"f3",x"49"),
  2247 => (x"c7",x"02",x"66",x"d4"),
  2248 => (x"87",x"da",x"49",x"87"),
  2249 => (x"87",x"c2",x"4a",x"70"),
  2250 => (x"cc",x"c2",x"4a",x"c0"),
  2251 => (x"f2",x"26",x"5a",x"fe"),
  2252 => (x"00",x"00",x"87",x"d9"),
  2253 => (x"00",x"00",x"00",x"00"),
  2254 => (x"00",x"00",x"00",x"00"),
  2255 => (x"71",x"1e",x"00",x"00"),
  2256 => (x"bf",x"c8",x"ff",x"4a"),
  2257 => (x"48",x"a1",x"72",x"49"),
  2258 => (x"ff",x"1e",x"4f",x"26"),
  2259 => (x"fe",x"89",x"bf",x"c8"),
  2260 => (x"c0",x"c0",x"c0",x"c0"),
  2261 => (x"c4",x"01",x"a9",x"c0"),
  2262 => (x"c2",x"4a",x"c0",x"87"),
  2263 => (x"72",x"4a",x"c1",x"87"),
  2264 => (x"1e",x"4f",x"26",x"48"),
  2265 => (x"bf",x"cc",x"ce",x"c2"),
  2266 => (x"c2",x"b9",x"c1",x"49"),
  2267 => (x"ff",x"59",x"d0",x"ce"),
  2268 => (x"ff",x"c3",x"48",x"d4"),
  2269 => (x"48",x"d0",x"ff",x"78"),
  2270 => (x"ff",x"78",x"e1",x"c0"),
  2271 => (x"78",x"c1",x"48",x"d4"),
  2272 => (x"78",x"71",x"31",x"c4"),
  2273 => (x"c0",x"48",x"d0",x"ff"),
  2274 => (x"4f",x"26",x"78",x"e0"),
  2275 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

