library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c4f2c287",
    12 => x"86c0c84e",
    13 => x"49c4f2c2",
    14 => x"48ccdfc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087d9e2",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"c44a711e",
    47 => x"c1484966",
    48 => x"58a6c888",
    49 => x"d4029971",
    50 => x"ff481287",
    51 => x"c47808d4",
    52 => x"c1484966",
    53 => x"58a6c888",
    54 => x"ec059971",
    55 => x"1e4f2687",
    56 => x"66c44a71",
    57 => x"88c14849",
    58 => x"7158a6c8",
    59 => x"87d60299",
    60 => x"c348d4ff",
    61 => x"526878ff",
    62 => x"484966c4",
    63 => x"a6c888c1",
    64 => x"05997158",
    65 => x"4f2687ea",
    66 => x"ff1e731e",
    67 => x"ffc34bd4",
    68 => x"c34a6b7b",
    69 => x"496b7bff",
    70 => x"b17232c8",
    71 => x"6b7bffc3",
    72 => x"7131c84a",
    73 => x"7bffc3b2",
    74 => x"32c8496b",
    75 => x"4871b172",
    76 => x"4d2687c4",
    77 => x"4b264c26",
    78 => x"5e0e4f26",
    79 => x"0e5d5c5b",
    80 => x"d4ff4a71",
    81 => x"c349724c",
    82 => x"7c7199ff",
    83 => x"bfccdfc2",
    84 => x"d087c805",
    85 => x"30c94866",
    86 => x"d058a6d4",
    87 => x"29d84966",
    88 => x"7199ffc3",
    89 => x"4966d07c",
    90 => x"ffc329d0",
    91 => x"d07c7199",
    92 => x"29c84966",
    93 => x"7199ffc3",
    94 => x"4966d07c",
    95 => x"7199ffc3",
    96 => x"d049727c",
    97 => x"99ffc329",
    98 => x"4b6c7c71",
    99 => x"4dfff0c9",
   100 => x"05abffc3",
   101 => x"ffc387d0",
   102 => x"c14b6c7c",
   103 => x"87c6028d",
   104 => x"02abffc3",
   105 => x"487387f0",
   106 => x"1e87c7fe",
   107 => x"d4ff49c0",
   108 => x"78ffc348",
   109 => x"c8c381c1",
   110 => x"f104a9b7",
   111 => x"1e4f2687",
   112 => x"87e71e73",
   113 => x"4bdff8c4",
   114 => x"ffc01ec0",
   115 => x"49f7c1f0",
   116 => x"c487e7fd",
   117 => x"05a8c186",
   118 => x"ff87eac0",
   119 => x"ffc348d4",
   120 => x"c0c0c178",
   121 => x"1ec0c0c0",
   122 => x"c1f0e1c0",
   123 => x"c9fd49e9",
   124 => x"7086c487",
   125 => x"87ca0598",
   126 => x"c348d4ff",
   127 => x"48c178ff",
   128 => x"e6fe87cb",
   129 => x"058bc187",
   130 => x"c087fdfe",
   131 => x"87e6fc48",
   132 => x"ff1e731e",
   133 => x"ffc348d4",
   134 => x"c04bd378",
   135 => x"f0ffc01e",
   136 => x"fc49c1c1",
   137 => x"86c487d4",
   138 => x"ca059870",
   139 => x"48d4ff87",
   140 => x"c178ffc3",
   141 => x"fd87cb48",
   142 => x"8bc187f1",
   143 => x"87dbff05",
   144 => x"f1fb48c0",
   145 => x"5b5e0e87",
   146 => x"d4ff0e5c",
   147 => x"87dbfd4c",
   148 => x"c01eeac6",
   149 => x"c8c1f0e1",
   150 => x"87defb49",
   151 => x"a8c186c4",
   152 => x"fe87c802",
   153 => x"48c087ea",
   154 => x"fa87e2c1",
   155 => x"497087da",
   156 => x"99ffffcf",
   157 => x"02a9eac6",
   158 => x"d3fe87c8",
   159 => x"c148c087",
   160 => x"ffc387cb",
   161 => x"4bf1c07c",
   162 => x"7087f4fc",
   163 => x"ebc00298",
   164 => x"c01ec087",
   165 => x"fac1f0ff",
   166 => x"87defa49",
   167 => x"987086c4",
   168 => x"c387d905",
   169 => x"496c7cff",
   170 => x"7c7cffc3",
   171 => x"c0c17c7c",
   172 => x"87c40299",
   173 => x"87d548c1",
   174 => x"87d148c0",
   175 => x"c405abc2",
   176 => x"c848c087",
   177 => x"058bc187",
   178 => x"c087fdfe",
   179 => x"87e4f948",
   180 => x"c21e731e",
   181 => x"c148ccdf",
   182 => x"ff4bc778",
   183 => x"78c248d0",
   184 => x"ff87c8fb",
   185 => x"78c348d0",
   186 => x"e5c01ec0",
   187 => x"49c0c1d0",
   188 => x"c487c7f9",
   189 => x"05a8c186",
   190 => x"c24b87c1",
   191 => x"87c505ab",
   192 => x"f9c048c0",
   193 => x"058bc187",
   194 => x"fc87d0ff",
   195 => x"dfc287f7",
   196 => x"987058d0",
   197 => x"c187cd05",
   198 => x"f0ffc01e",
   199 => x"f849d0c1",
   200 => x"86c487d8",
   201 => x"c348d4ff",
   202 => x"dec478ff",
   203 => x"d4dfc287",
   204 => x"48d0ff58",
   205 => x"d4ff78c2",
   206 => x"78ffc348",
   207 => x"f5f748c1",
   208 => x"5b5e0e87",
   209 => x"710e5d5c",
   210 => x"4dffc34a",
   211 => x"754cd4ff",
   212 => x"48d0ff7c",
   213 => x"7578c3c4",
   214 => x"c01e727c",
   215 => x"d8c1f0ff",
   216 => x"87d6f749",
   217 => x"987086c4",
   218 => x"c187c502",
   219 => x"87f0c048",
   220 => x"fec37c75",
   221 => x"1ec0c87c",
   222 => x"f44966d4",
   223 => x"86c487fa",
   224 => x"7c757c75",
   225 => x"dad87c75",
   226 => x"7c754be0",
   227 => x"0599496c",
   228 => x"8bc187c5",
   229 => x"7587f305",
   230 => x"48d0ff7c",
   231 => x"48c078c2",
   232 => x"0e87cff6",
   233 => x"5d5c5b5e",
   234 => x"c04b710e",
   235 => x"cdeec54c",
   236 => x"d4ff4adf",
   237 => x"78ffc348",
   238 => x"fec34968",
   239 => x"fdc005a9",
   240 => x"734d7087",
   241 => x"87cc029b",
   242 => x"731e66d0",
   243 => x"87cff449",
   244 => x"87d686c4",
   245 => x"c448d0ff",
   246 => x"ffc378d1",
   247 => x"4866d07d",
   248 => x"a6d488c1",
   249 => x"05987058",
   250 => x"d4ff87f0",
   251 => x"78ffc348",
   252 => x"059b7378",
   253 => x"d0ff87c5",
   254 => x"c178d048",
   255 => x"8ac14c4a",
   256 => x"87eefe05",
   257 => x"e9f44874",
   258 => x"1e731e87",
   259 => x"4bc04a71",
   260 => x"c348d4ff",
   261 => x"d0ff78ff",
   262 => x"78c3c448",
   263 => x"c348d4ff",
   264 => x"1e7278ff",
   265 => x"c1f0ffc0",
   266 => x"cdf449d1",
   267 => x"7086c487",
   268 => x"87d20598",
   269 => x"cc1ec0c8",
   270 => x"e6fd4966",
   271 => x"7086c487",
   272 => x"48d0ff4b",
   273 => x"487378c2",
   274 => x"0e87ebf3",
   275 => x"5d5c5b5e",
   276 => x"c01ec00e",
   277 => x"c9c1f0ff",
   278 => x"87def349",
   279 => x"dfc21ed2",
   280 => x"fefc49d4",
   281 => x"c086c887",
   282 => x"d284c14c",
   283 => x"f804acb7",
   284 => x"d4dfc287",
   285 => x"c349bf97",
   286 => x"c0c199c0",
   287 => x"e7c005a9",
   288 => x"dbdfc287",
   289 => x"d049bf97",
   290 => x"dcdfc231",
   291 => x"c84abf97",
   292 => x"c2b17232",
   293 => x"bf97dddf",
   294 => x"4c71b14a",
   295 => x"ffffffcf",
   296 => x"ca84c19c",
   297 => x"87e7c134",
   298 => x"97dddfc2",
   299 => x"31c149bf",
   300 => x"dfc299c6",
   301 => x"4abf97de",
   302 => x"722ab7c7",
   303 => x"d9dfc2b1",
   304 => x"4d4abf97",
   305 => x"dfc29dcf",
   306 => x"4abf97da",
   307 => x"32ca9ac3",
   308 => x"97dbdfc2",
   309 => x"33c24bbf",
   310 => x"dfc2b273",
   311 => x"4bbf97dc",
   312 => x"c69bc0c3",
   313 => x"b2732bb7",
   314 => x"48c181c2",
   315 => x"49703071",
   316 => x"307548c1",
   317 => x"4c724d70",
   318 => x"947184c1",
   319 => x"adb7c0c8",
   320 => x"c187cc06",
   321 => x"c82db734",
   322 => x"01adb7c0",
   323 => x"7487f4ff",
   324 => x"87def048",
   325 => x"5c5b5e0e",
   326 => x"86f80e5d",
   327 => x"48fae7c2",
   328 => x"dfc278c0",
   329 => x"49c01ef2",
   330 => x"c487defb",
   331 => x"05987086",
   332 => x"48c087c5",
   333 => x"c087cec9",
   334 => x"c07ec14d",
   335 => x"49bff6f2",
   336 => x"4ae8e0c2",
   337 => x"ec4bc871",
   338 => x"987087e0",
   339 => x"c087c205",
   340 => x"f2f2c07e",
   341 => x"e1c249bf",
   342 => x"c8714ac4",
   343 => x"87caec4b",
   344 => x"c2059870",
   345 => x"6e7ec087",
   346 => x"87fdc002",
   347 => x"bff8e6c2",
   348 => x"f0e7c24d",
   349 => x"487ebf9f",
   350 => x"a8ead6c5",
   351 => x"c287c705",
   352 => x"4dbff8e6",
   353 => x"486e87ce",
   354 => x"a8d5e9ca",
   355 => x"c087c502",
   356 => x"87f1c748",
   357 => x"1ef2dfc2",
   358 => x"ecf94975",
   359 => x"7086c487",
   360 => x"87c50598",
   361 => x"dcc748c0",
   362 => x"f2f2c087",
   363 => x"e1c249bf",
   364 => x"c8714ac4",
   365 => x"87f2ea4b",
   366 => x"c8059870",
   367 => x"fae7c287",
   368 => x"da78c148",
   369 => x"f6f2c087",
   370 => x"e0c249bf",
   371 => x"c8714ae8",
   372 => x"87d6ea4b",
   373 => x"c0029870",
   374 => x"48c087c5",
   375 => x"c287e6c6",
   376 => x"bf97f0e7",
   377 => x"a9d5c149",
   378 => x"87cdc005",
   379 => x"97f1e7c2",
   380 => x"eac249bf",
   381 => x"c5c002a9",
   382 => x"c648c087",
   383 => x"dfc287c7",
   384 => x"7ebf97f2",
   385 => x"a8e9c348",
   386 => x"87cec002",
   387 => x"ebc3486e",
   388 => x"c5c002a8",
   389 => x"c548c087",
   390 => x"dfc287eb",
   391 => x"49bf97fd",
   392 => x"ccc00599",
   393 => x"fedfc287",
   394 => x"c249bf97",
   395 => x"c5c002a9",
   396 => x"c548c087",
   397 => x"dfc287cf",
   398 => x"48bf97ff",
   399 => x"58f6e7c2",
   400 => x"c1484c70",
   401 => x"fae7c288",
   402 => x"c0e0c258",
   403 => x"7549bf97",
   404 => x"c1e0c281",
   405 => x"c84abf97",
   406 => x"7ea17232",
   407 => x"48c7ecc2",
   408 => x"e0c2786e",
   409 => x"48bf97c2",
   410 => x"c258a6c8",
   411 => x"02bffae7",
   412 => x"c087d4c2",
   413 => x"49bff2f2",
   414 => x"4ac4e1c2",
   415 => x"e74bc871",
   416 => x"987087e8",
   417 => x"87c5c002",
   418 => x"f8c348c0",
   419 => x"f2e7c287",
   420 => x"ecc24cbf",
   421 => x"e0c25cdb",
   422 => x"49bf97d7",
   423 => x"e0c231c8",
   424 => x"4abf97d6",
   425 => x"e0c249a1",
   426 => x"4abf97d8",
   427 => x"a17232d0",
   428 => x"d9e0c249",
   429 => x"d84abf97",
   430 => x"49a17232",
   431 => x"c29166c4",
   432 => x"81bfc7ec",
   433 => x"59cfecc2",
   434 => x"97dfe0c2",
   435 => x"32c84abf",
   436 => x"97dee0c2",
   437 => x"4aa24bbf",
   438 => x"97e0e0c2",
   439 => x"33d04bbf",
   440 => x"c24aa273",
   441 => x"bf97e1e0",
   442 => x"d89bcf4b",
   443 => x"4aa27333",
   444 => x"5ad3ecc2",
   445 => x"bfcfecc2",
   446 => x"748ac24a",
   447 => x"d3ecc292",
   448 => x"78a17248",
   449 => x"c287cac1",
   450 => x"bf97c4e0",
   451 => x"c231c849",
   452 => x"bf97c3e0",
   453 => x"c249a14a",
   454 => x"c259c2e8",
   455 => x"49bffee7",
   456 => x"ffc731c5",
   457 => x"c229c981",
   458 => x"c259dbec",
   459 => x"bf97c9e0",
   460 => x"c232c84a",
   461 => x"bf97c8e0",
   462 => x"c44aa24b",
   463 => x"826e9266",
   464 => x"5ad7ecc2",
   465 => x"48cfecc2",
   466 => x"ecc278c0",
   467 => x"a17248cb",
   468 => x"dbecc278",
   469 => x"cfecc248",
   470 => x"ecc278bf",
   471 => x"ecc248df",
   472 => x"c278bfd3",
   473 => x"02bffae7",
   474 => x"7487c9c0",
   475 => x"7030c448",
   476 => x"87c9c07e",
   477 => x"bfd7ecc2",
   478 => x"7030c448",
   479 => x"fee7c27e",
   480 => x"c1786e48",
   481 => x"268ef848",
   482 => x"264c264d",
   483 => x"0e4f264b",
   484 => x"5d5c5b5e",
   485 => x"c24a710e",
   486 => x"02bffae7",
   487 => x"4b7287cb",
   488 => x"4c722bc7",
   489 => x"c99cffc1",
   490 => x"c84b7287",
   491 => x"c34c722b",
   492 => x"ecc29cff",
   493 => x"c083bfc7",
   494 => x"abbfeef2",
   495 => x"c087d902",
   496 => x"c25bf2f2",
   497 => x"731ef2df",
   498 => x"87fdf049",
   499 => x"987086c4",
   500 => x"c087c505",
   501 => x"87e6c048",
   502 => x"bffae7c2",
   503 => x"7487d202",
   504 => x"c291c449",
   505 => x"6981f2df",
   506 => x"ffffcf4d",
   507 => x"cb9dffff",
   508 => x"c2497487",
   509 => x"f2dfc291",
   510 => x"4d699f81",
   511 => x"c6fe4875",
   512 => x"5b5e0e87",
   513 => x"f80e5d5c",
   514 => x"9c4c7186",
   515 => x"c087c505",
   516 => x"87c1c348",
   517 => x"6e7ea4c8",
   518 => x"d878c048",
   519 => x"87c70266",
   520 => x"bf9766d8",
   521 => x"c087c505",
   522 => x"87e9c248",
   523 => x"49c11ec0",
   524 => x"c487e0ca",
   525 => x"9d4d7086",
   526 => x"87c2c102",
   527 => x"4ac2e8c2",
   528 => x"e04966d8",
   529 => x"987087c9",
   530 => x"87f2c002",
   531 => x"66d84a75",
   532 => x"e04bcb49",
   533 => x"987087ee",
   534 => x"87e2c002",
   535 => x"9d751ec0",
   536 => x"c887c702",
   537 => x"78c048a6",
   538 => x"a6c887c5",
   539 => x"c878c148",
   540 => x"dec94966",
   541 => x"7086c487",
   542 => x"fe059d4d",
   543 => x"9d7587fe",
   544 => x"87cfc102",
   545 => x"6e49a5dc",
   546 => x"da786948",
   547 => x"a6c449a5",
   548 => x"78a4c448",
   549 => x"c448699f",
   550 => x"c2780866",
   551 => x"02bffae7",
   552 => x"a5d487d2",
   553 => x"49699f49",
   554 => x"99ffffc0",
   555 => x"30d04871",
   556 => x"87c27e70",
   557 => x"496e7ec0",
   558 => x"bf66c448",
   559 => x"0866c480",
   560 => x"cc7cc078",
   561 => x"66c449a4",
   562 => x"a4d079bf",
   563 => x"c179c049",
   564 => x"c087c248",
   565 => x"fa8ef848",
   566 => x"5e0e87ed",
   567 => x"0e5d5c5b",
   568 => x"029c4c71",
   569 => x"c887cac1",
   570 => x"026949a4",
   571 => x"d087c2c1",
   572 => x"496c4a66",
   573 => x"5aa6d482",
   574 => x"b94d66d0",
   575 => x"bff6e7c2",
   576 => x"72baff4a",
   577 => x"02997199",
   578 => x"c487e4c0",
   579 => x"496b4ba4",
   580 => x"7087fcf9",
   581 => x"f2e7c27b",
   582 => x"816c49bf",
   583 => x"b9757c71",
   584 => x"bff6e7c2",
   585 => x"72baff4a",
   586 => x"05997199",
   587 => x"7587dcff",
   588 => x"87d3f97c",
   589 => x"711e731e",
   590 => x"c7029b4b",
   591 => x"49a3c887",
   592 => x"87c50569",
   593 => x"f7c048c0",
   594 => x"cbecc287",
   595 => x"a3c44abf",
   596 => x"c2496949",
   597 => x"f2e7c289",
   598 => x"a27191bf",
   599 => x"f6e7c24a",
   600 => x"996b49bf",
   601 => x"c04aa271",
   602 => x"c85af2f2",
   603 => x"49721e66",
   604 => x"c487d6ea",
   605 => x"05987086",
   606 => x"48c087c4",
   607 => x"48c187c2",
   608 => x"1e87c8f8",
   609 => x"4b711e73",
   610 => x"87c7029b",
   611 => x"6949a3c8",
   612 => x"c087c505",
   613 => x"87f7c048",
   614 => x"bfcbecc2",
   615 => x"49a3c44a",
   616 => x"89c24969",
   617 => x"bff2e7c2",
   618 => x"4aa27191",
   619 => x"bff6e7c2",
   620 => x"71996b49",
   621 => x"f2c04aa2",
   622 => x"66c85af2",
   623 => x"e549721e",
   624 => x"86c487ff",
   625 => x"c4059870",
   626 => x"c248c087",
   627 => x"f648c187",
   628 => x"5e0e87f9",
   629 => x"1e0e5c5b",
   630 => x"66d04b71",
   631 => x"732cc94c",
   632 => x"d4c1029b",
   633 => x"49a3c887",
   634 => x"ccc10269",
   635 => x"f6e7c287",
   636 => x"b9ff49bf",
   637 => x"7e994a6b",
   638 => x"d103ac71",
   639 => x"d07bc087",
   640 => x"79c049a3",
   641 => x"c44aa3cc",
   642 => x"796a49a3",
   643 => x"8c7287c2",
   644 => x"c0029c74",
   645 => x"1e4987e3",
   646 => x"fdfa4973",
   647 => x"d086c487",
   648 => x"ffc74966",
   649 => x"87cb0299",
   650 => x"1ef2dfc2",
   651 => x"c3fc4973",
   652 => x"d086c487",
   653 => x"66d049a3",
   654 => x"ccf52679",
   655 => x"1e731e87",
   656 => x"029b4b71",
   657 => x"c287e4c0",
   658 => x"735bdfec",
   659 => x"c28ac24a",
   660 => x"49bff2e7",
   661 => x"cbecc292",
   662 => x"807248bf",
   663 => x"58e3ecc2",
   664 => x"30c44871",
   665 => x"58c2e8c2",
   666 => x"c287edc0",
   667 => x"c248dbec",
   668 => x"78bfcfec",
   669 => x"48dfecc2",
   670 => x"bfd3ecc2",
   671 => x"fae7c278",
   672 => x"87c902bf",
   673 => x"bff2e7c2",
   674 => x"c731c449",
   675 => x"d7ecc287",
   676 => x"31c449bf",
   677 => x"59c2e8c2",
   678 => x"0e87f0f3",
   679 => x"0e5c5b5e",
   680 => x"4bc04a71",
   681 => x"c0029a72",
   682 => x"a2da87e1",
   683 => x"4b699f49",
   684 => x"bffae7c2",
   685 => x"d487cf02",
   686 => x"699f49a2",
   687 => x"ffc04c49",
   688 => x"34d09cff",
   689 => x"4cc087c2",
   690 => x"73b34974",
   691 => x"87edfd49",
   692 => x"0e87f6f2",
   693 => x"5d5c5b5e",
   694 => x"7186f40e",
   695 => x"727ec04a",
   696 => x"87d8029a",
   697 => x"48eedfc2",
   698 => x"dfc278c0",
   699 => x"ecc248e6",
   700 => x"c278bfdf",
   701 => x"c248eadf",
   702 => x"78bfdbec",
   703 => x"48cfe8c2",
   704 => x"e7c250c0",
   705 => x"c249bffe",
   706 => x"4abfeedf",
   707 => x"c403aa71",
   708 => x"497287c9",
   709 => x"c00599cf",
   710 => x"f2c087e9",
   711 => x"dfc248ee",
   712 => x"c278bfe6",
   713 => x"c21ef2df",
   714 => x"49bfe6df",
   715 => x"48e6dfc2",
   716 => x"7178a1c1",
   717 => x"c487d2e3",
   718 => x"eaf2c086",
   719 => x"f2dfc248",
   720 => x"c087cc78",
   721 => x"48bfeaf2",
   722 => x"c080e0c0",
   723 => x"c258eef2",
   724 => x"48bfeedf",
   725 => x"dfc280c1",
   726 => x"aa2758f2",
   727 => x"bf00000c",
   728 => x"9d4dbf97",
   729 => x"87e3c202",
   730 => x"02ade5c3",
   731 => x"c087dcc2",
   732 => x"4bbfeaf2",
   733 => x"1149a3cb",
   734 => x"05accf4c",
   735 => x"7587d2c1",
   736 => x"c199df49",
   737 => x"c291cd89",
   738 => x"c181c2e8",
   739 => x"51124aa3",
   740 => x"124aa3c3",
   741 => x"4aa3c551",
   742 => x"a3c75112",
   743 => x"c951124a",
   744 => x"51124aa3",
   745 => x"124aa3ce",
   746 => x"4aa3d051",
   747 => x"a3d25112",
   748 => x"d451124a",
   749 => x"51124aa3",
   750 => x"124aa3d6",
   751 => x"4aa3d851",
   752 => x"a3dc5112",
   753 => x"de51124a",
   754 => x"51124aa3",
   755 => x"fac07ec1",
   756 => x"c8497487",
   757 => x"ebc00599",
   758 => x"d0497487",
   759 => x"87d10599",
   760 => x"c00266dc",
   761 => x"497387cb",
   762 => x"700f66dc",
   763 => x"d3c00298",
   764 => x"c0056e87",
   765 => x"e8c287c6",
   766 => x"50c048c2",
   767 => x"bfeaf2c0",
   768 => x"87e1c248",
   769 => x"48cfe8c2",
   770 => x"c27e50c0",
   771 => x"49bffee7",
   772 => x"bfeedfc2",
   773 => x"04aa714a",
   774 => x"c287f7fb",
   775 => x"05bfdfec",
   776 => x"c287c8c0",
   777 => x"02bffae7",
   778 => x"c287f8c1",
   779 => x"49bfeadf",
   780 => x"7087dced",
   781 => x"eedfc249",
   782 => x"48a6c459",
   783 => x"bfeadfc2",
   784 => x"fae7c278",
   785 => x"d8c002bf",
   786 => x"4966c487",
   787 => x"ffffffcf",
   788 => x"02a999f8",
   789 => x"c087c5c0",
   790 => x"87e1c04c",
   791 => x"dcc04cc1",
   792 => x"4966c487",
   793 => x"99f8ffcf",
   794 => x"c8c002a9",
   795 => x"48a6c887",
   796 => x"c5c078c0",
   797 => x"48a6c887",
   798 => x"66c878c1",
   799 => x"059c744c",
   800 => x"c487e0c0",
   801 => x"89c24966",
   802 => x"bff2e7c2",
   803 => x"ecc2914a",
   804 => x"c24abfcb",
   805 => x"7248e6df",
   806 => x"dfc278a1",
   807 => x"78c048ee",
   808 => x"c087dff9",
   809 => x"eb8ef448",
   810 => x"000087dd",
   811 => x"ffff0000",
   812 => x"0cbaffff",
   813 => x"0cc30000",
   814 => x"41460000",
   815 => x"20323354",
   816 => x"46002020",
   817 => x"36315441",
   818 => x"00202020",
   819 => x"48d4ff1e",
   820 => x"6878ffc3",
   821 => x"1e4f2648",
   822 => x"c348d4ff",
   823 => x"d0ff78ff",
   824 => x"78e1c048",
   825 => x"d448d4ff",
   826 => x"e3ecc278",
   827 => x"bfd4ff48",
   828 => x"1e4f2650",
   829 => x"c048d0ff",
   830 => x"4f2678e0",
   831 => x"87ccff1e",
   832 => x"02994970",
   833 => x"fbc087c6",
   834 => x"87f105a9",
   835 => x"4f264871",
   836 => x"5c5b5e0e",
   837 => x"c04b710e",
   838 => x"87f0fe4c",
   839 => x"02994970",
   840 => x"c087f9c0",
   841 => x"c002a9ec",
   842 => x"fbc087f2",
   843 => x"ebc002a9",
   844 => x"b766cc87",
   845 => x"87c703ac",
   846 => x"c20266d0",
   847 => x"71537187",
   848 => x"87c20299",
   849 => x"c3fe84c1",
   850 => x"99497087",
   851 => x"c087cd02",
   852 => x"c702a9ec",
   853 => x"a9fbc087",
   854 => x"87d5ff05",
   855 => x"c30266d0",
   856 => x"7b97c087",
   857 => x"05a9ecc0",
   858 => x"4a7487c4",
   859 => x"4a7487c5",
   860 => x"728a0ac0",
   861 => x"2687c248",
   862 => x"264c264d",
   863 => x"1e4f264b",
   864 => x"7087c9fd",
   865 => x"f0c04a49",
   866 => x"87c904aa",
   867 => x"01aaf9c0",
   868 => x"f0c087c3",
   869 => x"aac1c18a",
   870 => x"c187c904",
   871 => x"c301aada",
   872 => x"8af7c087",
   873 => x"04aae1c1",
   874 => x"fac187c9",
   875 => x"87c301aa",
   876 => x"728afdc0",
   877 => x"0e4f2648",
   878 => x"0e5c5b5e",
   879 => x"d4ff4a71",
   880 => x"c049724c",
   881 => x"4b7087e9",
   882 => x"87c2029b",
   883 => x"d0ff8bc1",
   884 => x"c178c548",
   885 => x"49737cd5",
   886 => x"e3c131c6",
   887 => x"4abf97fa",
   888 => x"70b07148",
   889 => x"48d0ff7c",
   890 => x"487378c4",
   891 => x"0e87cafe",
   892 => x"5d5c5b5e",
   893 => x"7186f80e",
   894 => x"fb7ec04c",
   895 => x"4bc087d9",
   896 => x"97dcfac0",
   897 => x"a9c049bf",
   898 => x"fb87cf04",
   899 => x"83c187ee",
   900 => x"97dcfac0",
   901 => x"06ab49bf",
   902 => x"fac087f1",
   903 => x"02bf97dc",
   904 => x"e7fa87cf",
   905 => x"99497087",
   906 => x"c087c602",
   907 => x"f105a9ec",
   908 => x"fa4bc087",
   909 => x"4d7087d6",
   910 => x"c887d1fa",
   911 => x"cbfa58a6",
   912 => x"c14a7087",
   913 => x"49a4c883",
   914 => x"ad496997",
   915 => x"c087c702",
   916 => x"c005adff",
   917 => x"a4c987e7",
   918 => x"49699749",
   919 => x"02a966c4",
   920 => x"c04887c7",
   921 => x"d405a8ff",
   922 => x"49a4ca87",
   923 => x"aa496997",
   924 => x"c087c602",
   925 => x"c405aaff",
   926 => x"d07ec187",
   927 => x"adecc087",
   928 => x"c087c602",
   929 => x"c405adfb",
   930 => x"c14bc087",
   931 => x"fe026e7e",
   932 => x"def987e1",
   933 => x"f8487387",
   934 => x"87dbfb8e",
   935 => x"5b5e0e00",
   936 => x"f80e5d5c",
   937 => x"ff4d7186",
   938 => x"1e754bd4",
   939 => x"49e8ecc2",
   940 => x"c487cee5",
   941 => x"02987086",
   942 => x"c487ccc4",
   943 => x"e3c148a6",
   944 => x"7578bffc",
   945 => x"87effb49",
   946 => x"c548d0ff",
   947 => x"7bd6c178",
   948 => x"a2754ac0",
   949 => x"c17b1149",
   950 => x"aab7cb82",
   951 => x"cc87f304",
   952 => x"7bffc34a",
   953 => x"e0c082c1",
   954 => x"f404aab7",
   955 => x"48d0ff87",
   956 => x"ffc378c4",
   957 => x"c178c57b",
   958 => x"7bc17bd3",
   959 => x"486678c4",
   960 => x"06a8b7c0",
   961 => x"c287f0c2",
   962 => x"4cbff0ec",
   963 => x"744866c4",
   964 => x"58a6c888",
   965 => x"c1029c74",
   966 => x"dfc287f9",
   967 => x"c0c87ef2",
   968 => x"b7c08c4d",
   969 => x"87c603ac",
   970 => x"4da4c0c8",
   971 => x"ecc24cc0",
   972 => x"49bf97e3",
   973 => x"d10299d0",
   974 => x"c21ec087",
   975 => x"e749e8ec",
   976 => x"86c487f2",
   977 => x"c04a4970",
   978 => x"dfc287ee",
   979 => x"ecc21ef2",
   980 => x"dfe749e8",
   981 => x"7086c487",
   982 => x"d0ff4a49",
   983 => x"78c5c848",
   984 => x"6e7bd4c1",
   985 => x"6e7bbf97",
   986 => x"7080c148",
   987 => x"058dc17e",
   988 => x"ff87f0ff",
   989 => x"78c448d0",
   990 => x"c5059a72",
   991 => x"c148c087",
   992 => x"1ec187c7",
   993 => x"49e8ecc2",
   994 => x"c487cfe5",
   995 => x"059c7486",
   996 => x"c487c7fe",
   997 => x"b7c04866",
   998 => x"87d106a8",
   999 => x"48e8ecc2",
  1000 => x"80d078c0",
  1001 => x"80f478c0",
  1002 => x"bff4ecc2",
  1003 => x"4866c478",
  1004 => x"01a8b7c0",
  1005 => x"ff87d0fd",
  1006 => x"78c548d0",
  1007 => x"c07bd3c1",
  1008 => x"c178c47b",
  1009 => x"c087c248",
  1010 => x"268ef848",
  1011 => x"264c264d",
  1012 => x"0e4f264b",
  1013 => x"5d5c5b5e",
  1014 => x"4b711e0e",
  1015 => x"ab4d4cc0",
  1016 => x"87e8c004",
  1017 => x"1eeff7c0",
  1018 => x"c4029d75",
  1019 => x"c24ac087",
  1020 => x"724ac187",
  1021 => x"87dbeb49",
  1022 => x"7e7086c4",
  1023 => x"056e84c1",
  1024 => x"4c7387c2",
  1025 => x"ac7385c1",
  1026 => x"87d8ff06",
  1027 => x"fe26486e",
  1028 => x"5e0e87f9",
  1029 => x"710e5c5b",
  1030 => x"0266cc4b",
  1031 => x"c04c87d8",
  1032 => x"d8028cf0",
  1033 => x"c14a7487",
  1034 => x"87d1028a",
  1035 => x"87cd028a",
  1036 => x"87c9028a",
  1037 => x"497387d9",
  1038 => x"d287e2f9",
  1039 => x"c01e7487",
  1040 => x"d9dbc149",
  1041 => x"731e7487",
  1042 => x"d1dbc149",
  1043 => x"fd86c887",
  1044 => x"5e0e87fb",
  1045 => x"0e5d5c5b",
  1046 => x"494c711e",
  1047 => x"edc291de",
  1048 => x"85714dd0",
  1049 => x"c1026d97",
  1050 => x"ecc287dc",
  1051 => x"744abffc",
  1052 => x"fd497282",
  1053 => x"7e7087dd",
  1054 => x"f2c0026e",
  1055 => x"c4edc287",
  1056 => x"cb4a6e4b",
  1057 => x"dfc0ff49",
  1058 => x"cb4b7487",
  1059 => x"cee4c193",
  1060 => x"c183c483",
  1061 => x"747bcac3",
  1062 => x"d1c5c149",
  1063 => x"c17b7587",
  1064 => x"bf97fbe3",
  1065 => x"edc21e49",
  1066 => x"e5fd49c4",
  1067 => x"7486c487",
  1068 => x"f9c4c149",
  1069 => x"c149c087",
  1070 => x"c287d8c6",
  1071 => x"c048e4ec",
  1072 => x"dd49c178",
  1073 => x"fc2687d9",
  1074 => x"6f4c87c1",
  1075 => x"6e696461",
  1076 => x"2e2e2e67",
  1077 => x"5b5e0e00",
  1078 => x"4b710e5c",
  1079 => x"fcecc24a",
  1080 => x"497282bf",
  1081 => x"7087ecfb",
  1082 => x"c4029c4c",
  1083 => x"eae64987",
  1084 => x"fcecc287",
  1085 => x"c178c048",
  1086 => x"87e3dc49",
  1087 => x"0e87cefb",
  1088 => x"5d5c5b5e",
  1089 => x"c286f40e",
  1090 => x"c04df2df",
  1091 => x"48a6c44c",
  1092 => x"ecc278c0",
  1093 => x"c049bffc",
  1094 => x"c1c106a9",
  1095 => x"f2dfc287",
  1096 => x"c0029848",
  1097 => x"f7c087f8",
  1098 => x"66c81eef",
  1099 => x"c487c702",
  1100 => x"78c048a6",
  1101 => x"a6c487c5",
  1102 => x"c478c148",
  1103 => x"d2e64966",
  1104 => x"7086c487",
  1105 => x"c484c14d",
  1106 => x"80c14866",
  1107 => x"c258a6c8",
  1108 => x"49bffcec",
  1109 => x"87c603ac",
  1110 => x"ff059d75",
  1111 => x"4cc087c8",
  1112 => x"c3029d75",
  1113 => x"f7c087e0",
  1114 => x"66c81eef",
  1115 => x"cc87c702",
  1116 => x"78c048a6",
  1117 => x"a6cc87c5",
  1118 => x"cc78c148",
  1119 => x"d2e54966",
  1120 => x"7086c487",
  1121 => x"c2026e7e",
  1122 => x"496e87e9",
  1123 => x"699781cb",
  1124 => x"0299d049",
  1125 => x"c187d6c1",
  1126 => x"744ad5c3",
  1127 => x"c191cb49",
  1128 => x"7281cee4",
  1129 => x"c381c879",
  1130 => x"497451ff",
  1131 => x"edc291de",
  1132 => x"85714dd0",
  1133 => x"7d97c1c2",
  1134 => x"c049a5c1",
  1135 => x"e8c251e0",
  1136 => x"02bf97c2",
  1137 => x"84c187d2",
  1138 => x"c24ba5c2",
  1139 => x"db4ac2e8",
  1140 => x"d3fbfe49",
  1141 => x"87dbc187",
  1142 => x"c049a5cd",
  1143 => x"c284c151",
  1144 => x"4a6e4ba5",
  1145 => x"fafe49cb",
  1146 => x"c6c187fe",
  1147 => x"d2c1c187",
  1148 => x"cb49744a",
  1149 => x"cee4c191",
  1150 => x"c2797281",
  1151 => x"bf97c2e8",
  1152 => x"7487d802",
  1153 => x"c191de49",
  1154 => x"d0edc284",
  1155 => x"c283714b",
  1156 => x"dd4ac2e8",
  1157 => x"cffafe49",
  1158 => x"7487d887",
  1159 => x"c293de4b",
  1160 => x"cb83d0ed",
  1161 => x"51c049a3",
  1162 => x"6e7384c1",
  1163 => x"fe49cb4a",
  1164 => x"c487f5f9",
  1165 => x"80c14866",
  1166 => x"c758a6c8",
  1167 => x"c5c003ac",
  1168 => x"fc056e87",
  1169 => x"487487e0",
  1170 => x"fef58ef4",
  1171 => x"1e731e87",
  1172 => x"cb494b71",
  1173 => x"cee4c191",
  1174 => x"4aa1c881",
  1175 => x"48fae3c1",
  1176 => x"a1c95012",
  1177 => x"dcfac04a",
  1178 => x"ca501248",
  1179 => x"fbe3c181",
  1180 => x"c1501148",
  1181 => x"bf97fbe3",
  1182 => x"49c01e49",
  1183 => x"c287d3f6",
  1184 => x"de48e4ec",
  1185 => x"d649c178",
  1186 => x"f52687d5",
  1187 => x"711e87c1",
  1188 => x"91cb494a",
  1189 => x"81cee4c1",
  1190 => x"481181c8",
  1191 => x"58e8ecc2",
  1192 => x"48fcecc2",
  1193 => x"49c178c0",
  1194 => x"2687f4d5",
  1195 => x"49c01e4f",
  1196 => x"87dffec0",
  1197 => x"711e4f26",
  1198 => x"87d20299",
  1199 => x"48e3e5c1",
  1200 => x"80f750c0",
  1201 => x"40cecac1",
  1202 => x"78c7e4c1",
  1203 => x"e5c187ce",
  1204 => x"e4c148df",
  1205 => x"80fc78c0",
  1206 => x"78edcac1",
  1207 => x"5e0e4f26",
  1208 => x"710e5c5b",
  1209 => x"92cb4a4c",
  1210 => x"82cee4c1",
  1211 => x"c949a2c8",
  1212 => x"6b974ba2",
  1213 => x"69971e4b",
  1214 => x"82ca1e49",
  1215 => x"e7c04912",
  1216 => x"49c087d8",
  1217 => x"7487d8d4",
  1218 => x"e1fbc049",
  1219 => x"f28ef887",
  1220 => x"731e87fb",
  1221 => x"494b711e",
  1222 => x"7387c3ff",
  1223 => x"87fefe49",
  1224 => x"1e87ecf2",
  1225 => x"4b711e73",
  1226 => x"024aa3c6",
  1227 => x"8ac187db",
  1228 => x"8a87d602",
  1229 => x"87dac102",
  1230 => x"fcc0028a",
  1231 => x"c0028a87",
  1232 => x"028a87e1",
  1233 => x"dbc187cb",
  1234 => x"fd49c787",
  1235 => x"dec187c0",
  1236 => x"fcecc287",
  1237 => x"cbc102bf",
  1238 => x"88c14887",
  1239 => x"58c0edc2",
  1240 => x"c287c1c1",
  1241 => x"02bfc0ed",
  1242 => x"c287f9c0",
  1243 => x"48bffcec",
  1244 => x"edc280c1",
  1245 => x"ebc058c0",
  1246 => x"fcecc287",
  1247 => x"89c649bf",
  1248 => x"59c0edc2",
  1249 => x"03a9b7c0",
  1250 => x"ecc287da",
  1251 => x"78c048fc",
  1252 => x"edc287d2",
  1253 => x"cb02bfc0",
  1254 => x"fcecc287",
  1255 => x"80c648bf",
  1256 => x"58c0edc2",
  1257 => x"f6d149c0",
  1258 => x"c0497387",
  1259 => x"f087fff8",
  1260 => x"5e0e87dd",
  1261 => x"0e5d5c5b",
  1262 => x"dc86d0ff",
  1263 => x"a6c859a6",
  1264 => x"c478c048",
  1265 => x"66c4c180",
  1266 => x"c180c478",
  1267 => x"c180c478",
  1268 => x"c0edc278",
  1269 => x"c278c148",
  1270 => x"48bfe4ec",
  1271 => x"cb05a8de",
  1272 => x"87dbf487",
  1273 => x"a6cc4970",
  1274 => x"87f2cf59",
  1275 => x"e487e8e3",
  1276 => x"d7e387ca",
  1277 => x"c04c7087",
  1278 => x"c102acfb",
  1279 => x"66d887fb",
  1280 => x"87edc105",
  1281 => x"4a66c0c1",
  1282 => x"7e6a82c4",
  1283 => x"e0c11e72",
  1284 => x"66c448d3",
  1285 => x"4aa1c849",
  1286 => x"aa714120",
  1287 => x"1087f905",
  1288 => x"c14a2651",
  1289 => x"c14866c0",
  1290 => x"6a78cdc9",
  1291 => x"7481c749",
  1292 => x"66c0c151",
  1293 => x"c181c849",
  1294 => x"66c0c151",
  1295 => x"c081c949",
  1296 => x"66c0c151",
  1297 => x"c081ca49",
  1298 => x"d81ec151",
  1299 => x"c8496a1e",
  1300 => x"87fce281",
  1301 => x"c4c186c8",
  1302 => x"a8c04866",
  1303 => x"c887c701",
  1304 => x"78c148a6",
  1305 => x"c4c187ce",
  1306 => x"88c14866",
  1307 => x"c358a6d0",
  1308 => x"87c8e287",
  1309 => x"c248a6d0",
  1310 => x"029c7478",
  1311 => x"c887dbcd",
  1312 => x"c8c14866",
  1313 => x"cd03a866",
  1314 => x"a6dc87d0",
  1315 => x"e878c048",
  1316 => x"e078c080",
  1317 => x"4c7087f6",
  1318 => x"05acd0c1",
  1319 => x"c487d9c2",
  1320 => x"dae37e66",
  1321 => x"c8497087",
  1322 => x"dfe059a6",
  1323 => x"c04c7087",
  1324 => x"c105acec",
  1325 => x"66c887ed",
  1326 => x"c191cb49",
  1327 => x"c48166c0",
  1328 => x"4d6a4aa1",
  1329 => x"c44aa1c8",
  1330 => x"cac15266",
  1331 => x"dfff79ce",
  1332 => x"4c7087fa",
  1333 => x"87d9029c",
  1334 => x"02acfbc0",
  1335 => x"557487d3",
  1336 => x"87e8dfff",
  1337 => x"029c4c70",
  1338 => x"fbc087c7",
  1339 => x"edff05ac",
  1340 => x"55e0c087",
  1341 => x"c055c1c2",
  1342 => x"66d87d97",
  1343 => x"05a96e49",
  1344 => x"66c887db",
  1345 => x"a866cc48",
  1346 => x"c887ca04",
  1347 => x"80c14866",
  1348 => x"c858a6cc",
  1349 => x"4866cc87",
  1350 => x"a6d088c1",
  1351 => x"ebdeff58",
  1352 => x"c14c7087",
  1353 => x"c805acd0",
  1354 => x"4866d487",
  1355 => x"a6d880c1",
  1356 => x"acd0c158",
  1357 => x"87e7fd02",
  1358 => x"48a6e0c0",
  1359 => x"c47866d8",
  1360 => x"e0c04866",
  1361 => x"c905a866",
  1362 => x"e4c087e2",
  1363 => x"78c048a6",
  1364 => x"78c080c4",
  1365 => x"fbc04874",
  1366 => x"6e7e7088",
  1367 => x"87e5c802",
  1368 => x"88cb486e",
  1369 => x"026e7e70",
  1370 => x"6e87cdc1",
  1371 => x"7088c948",
  1372 => x"c3026e7e",
  1373 => x"486e87e9",
  1374 => x"7e7088c4",
  1375 => x"87ce026e",
  1376 => x"88c1486e",
  1377 => x"026e7e70",
  1378 => x"c787d4c3",
  1379 => x"a6dc87f1",
  1380 => x"78f0c048",
  1381 => x"87f4dcff",
  1382 => x"ecc04c70",
  1383 => x"c4c002ac",
  1384 => x"a6e0c087",
  1385 => x"acecc05c",
  1386 => x"ff87cd02",
  1387 => x"7087dddc",
  1388 => x"acecc04c",
  1389 => x"87f3ff05",
  1390 => x"02acecc0",
  1391 => x"ff87c4c0",
  1392 => x"c087c9dc",
  1393 => x"d01eca1e",
  1394 => x"91cb4966",
  1395 => x"4866c8c1",
  1396 => x"a6cc8071",
  1397 => x"4866c858",
  1398 => x"a6d080c4",
  1399 => x"bf66cc58",
  1400 => x"ebdcff49",
  1401 => x"de1ec187",
  1402 => x"bf66d41e",
  1403 => x"dfdcff49",
  1404 => x"7086d087",
  1405 => x"8909c049",
  1406 => x"59a6ecc0",
  1407 => x"4866e8c0",
  1408 => x"c006a8c0",
  1409 => x"e8c087ee",
  1410 => x"a8dd4866",
  1411 => x"87e4c003",
  1412 => x"49bf66c4",
  1413 => x"8166e8c0",
  1414 => x"c051e0c0",
  1415 => x"c14966e8",
  1416 => x"bf66c481",
  1417 => x"51c1c281",
  1418 => x"4966e8c0",
  1419 => x"66c481c2",
  1420 => x"51c081bf",
  1421 => x"c9c1486e",
  1422 => x"496e78cd",
  1423 => x"66d081c8",
  1424 => x"c9496e51",
  1425 => x"5166d481",
  1426 => x"81ca496e",
  1427 => x"d05166dc",
  1428 => x"80c14866",
  1429 => x"4858a6d4",
  1430 => x"78c180d8",
  1431 => x"ff87e6c4",
  1432 => x"7087dcdc",
  1433 => x"a6ecc049",
  1434 => x"d2dcff59",
  1435 => x"c0497087",
  1436 => x"dc59a6e0",
  1437 => x"ecc04866",
  1438 => x"cac005a8",
  1439 => x"48a6dc87",
  1440 => x"7866e8c0",
  1441 => x"ff87c4c0",
  1442 => x"c887c1d9",
  1443 => x"91cb4966",
  1444 => x"4866c0c1",
  1445 => x"7e708071",
  1446 => x"81c8496e",
  1447 => x"82ca4a6e",
  1448 => x"5266e8c0",
  1449 => x"c14a66dc",
  1450 => x"66e8c082",
  1451 => x"7248c18a",
  1452 => x"c14a7030",
  1453 => x"7997728a",
  1454 => x"1e496997",
  1455 => x"4966ecc0",
  1456 => x"c487d9d7",
  1457 => x"a6f0c086",
  1458 => x"c4496e58",
  1459 => x"c04d6981",
  1460 => x"c44866e0",
  1461 => x"c002a866",
  1462 => x"a6c487c8",
  1463 => x"c078c048",
  1464 => x"a6c487c5",
  1465 => x"c478c148",
  1466 => x"e0c01e66",
  1467 => x"ff49751e",
  1468 => x"c887ddd8",
  1469 => x"c04c7086",
  1470 => x"c106acb7",
  1471 => x"857487d4",
  1472 => x"7449e0c0",
  1473 => x"c14b7589",
  1474 => x"714adce0",
  1475 => x"87d8e6fe",
  1476 => x"e4c085c2",
  1477 => x"80c14866",
  1478 => x"58a6e8c0",
  1479 => x"4966ecc0",
  1480 => x"a97081c1",
  1481 => x"87c8c002",
  1482 => x"c048a6c4",
  1483 => x"87c5c078",
  1484 => x"c148a6c4",
  1485 => x"1e66c478",
  1486 => x"c049a4c2",
  1487 => x"887148e0",
  1488 => x"751e4970",
  1489 => x"c7d7ff49",
  1490 => x"c086c887",
  1491 => x"ff01a8b7",
  1492 => x"e4c087c0",
  1493 => x"d1c00266",
  1494 => x"c9496e87",
  1495 => x"66e4c081",
  1496 => x"c1486e51",
  1497 => x"c078decb",
  1498 => x"496e87cc",
  1499 => x"51c281c9",
  1500 => x"ccc1486e",
  1501 => x"e8c078d2",
  1502 => x"78c148a6",
  1503 => x"ff87c6c0",
  1504 => x"7087f9d5",
  1505 => x"66e8c04c",
  1506 => x"87f5c002",
  1507 => x"cc4866c8",
  1508 => x"c004a866",
  1509 => x"66c887cb",
  1510 => x"cc80c148",
  1511 => x"e0c058a6",
  1512 => x"4866cc87",
  1513 => x"a6d088c1",
  1514 => x"87d5c058",
  1515 => x"05acc6c1",
  1516 => x"d087c8c0",
  1517 => x"80c14866",
  1518 => x"ff58a6d4",
  1519 => x"7087fdd4",
  1520 => x"4866d44c",
  1521 => x"a6d880c1",
  1522 => x"029c7458",
  1523 => x"c887cbc0",
  1524 => x"c8c14866",
  1525 => x"f204a866",
  1526 => x"d4ff87f0",
  1527 => x"66c887d5",
  1528 => x"03a8c748",
  1529 => x"c287e5c0",
  1530 => x"c048c0ed",
  1531 => x"4966c878",
  1532 => x"c0c191cb",
  1533 => x"a1c48166",
  1534 => x"c04a6a4a",
  1535 => x"66c87952",
  1536 => x"cc80c148",
  1537 => x"a8c758a6",
  1538 => x"87dbff04",
  1539 => x"ff8ed0ff",
  1540 => x"4c87f8de",
  1541 => x"2064616f",
  1542 => x"00202e2a",
  1543 => x"1e00203a",
  1544 => x"4b711e73",
  1545 => x"87c6029b",
  1546 => x"48fcecc2",
  1547 => x"1ec778c0",
  1548 => x"bffcecc2",
  1549 => x"e4c11e49",
  1550 => x"ecc21ece",
  1551 => x"ed49bfe4",
  1552 => x"86cc87f0",
  1553 => x"bfe4ecc2",
  1554 => x"87eae949",
  1555 => x"c8029b73",
  1556 => x"cee4c187",
  1557 => x"e7e7c049",
  1558 => x"f2ddff87",
  1559 => x"e3c11e87",
  1560 => x"50c048fa",
  1561 => x"bff1e5c1",
  1562 => x"f0d8ff49",
  1563 => x"2648c087",
  1564 => x"e3c71e4f",
  1565 => x"fe49c187",
  1566 => x"e9fe87e5",
  1567 => x"987087d2",
  1568 => x"fe87cd02",
  1569 => x"7087cdf2",
  1570 => x"87c40298",
  1571 => x"87c24ac1",
  1572 => x"9a724ac0",
  1573 => x"c087ce05",
  1574 => x"c1e3c11e",
  1575 => x"f7f2c049",
  1576 => x"fe86c487",
  1577 => x"c11ec087",
  1578 => x"c049cce3",
  1579 => x"c087e9f2",
  1580 => x"87e9fe1e",
  1581 => x"f2c04970",
  1582 => x"dac387de",
  1583 => x"268ef887",
  1584 => x"2044534f",
  1585 => x"6c696166",
  1586 => x"002e6465",
  1587 => x"746f6f42",
  1588 => x"2e676e69",
  1589 => x"1e002e2e",
  1590 => x"87c0eac0",
  1591 => x"87eef5c0",
  1592 => x"4f2687f6",
  1593 => x"fcecc21e",
  1594 => x"c278c048",
  1595 => x"c048e4ec",
  1596 => x"87fdfd78",
  1597 => x"48c087e1",
  1598 => x"00004f26",
  1599 => x"00000001",
  1600 => x"78452080",
  1601 => x"80007469",
  1602 => x"63614220",
  1603 => x"128e006b",
  1604 => x"2b500000",
  1605 => x"00000000",
  1606 => x"00128e00",
  1607 => x"002b6e00",
  1608 => x"00000000",
  1609 => x"0000128e",
  1610 => x"00002b8c",
  1611 => x"8e000000",
  1612 => x"aa000012",
  1613 => x"0000002b",
  1614 => x"128e0000",
  1615 => x"2bc80000",
  1616 => x"00000000",
  1617 => x"00128e00",
  1618 => x"002be600",
  1619 => x"00000000",
  1620 => x"0000128e",
  1621 => x"00002c04",
  1622 => x"8e000000",
  1623 => x"00000012",
  1624 => x"00000000",
  1625 => x"13230000",
  1626 => x"00000000",
  1627 => x"00000000",
  1628 => x"00197500",
  1629 => x"34364300",
  1630 => x"20202020",
  1631 => x"4d4f5220",
  1632 => x"f0fe1e00",
  1633 => x"cd78c048",
  1634 => x"26097909",
  1635 => x"fe1e1e4f",
  1636 => x"487ebff0",
  1637 => x"1e4f2626",
  1638 => x"c148f0fe",
  1639 => x"1e4f2678",
  1640 => x"c048f0fe",
  1641 => x"1e4f2678",
  1642 => x"52c04a71",
  1643 => x"0e4f2652",
  1644 => x"5d5c5b5e",
  1645 => x"7186f40e",
  1646 => x"7e6d974d",
  1647 => x"974ca5c1",
  1648 => x"a6c8486c",
  1649 => x"c4486e58",
  1650 => x"c505a866",
  1651 => x"c048ff87",
  1652 => x"caff87e6",
  1653 => x"49a5c287",
  1654 => x"714b6c97",
  1655 => x"6b974ba3",
  1656 => x"7e6c974b",
  1657 => x"80c1486e",
  1658 => x"c758a6c8",
  1659 => x"58a6cc98",
  1660 => x"fe7c9770",
  1661 => x"487387e1",
  1662 => x"4d268ef4",
  1663 => x"4b264c26",
  1664 => x"5e0e4f26",
  1665 => x"f40e5c5b",
  1666 => x"d84c7186",
  1667 => x"ffc34a66",
  1668 => x"4ba4c29a",
  1669 => x"73496c97",
  1670 => x"517249a1",
  1671 => x"6e7e6c97",
  1672 => x"c880c148",
  1673 => x"98c758a6",
  1674 => x"7058a6cc",
  1675 => x"ff8ef454",
  1676 => x"1e1e87ca",
  1677 => x"e087e8fd",
  1678 => x"c0494abf",
  1679 => x"0299c0e0",
  1680 => x"1e7287cb",
  1681 => x"49e2f0c2",
  1682 => x"c487f7fe",
  1683 => x"87fdfc86",
  1684 => x"c2fd7e70",
  1685 => x"4f262687",
  1686 => x"e2f0c21e",
  1687 => x"87c7fd49",
  1688 => x"49f2e8c1",
  1689 => x"c487dafc",
  1690 => x"4f2687c7",
  1691 => x"48d0ff1e",
  1692 => x"ff78e1c8",
  1693 => x"78c548d4",
  1694 => x"c30266c4",
  1695 => x"78e0c387",
  1696 => x"c60266c8",
  1697 => x"48d4ff87",
  1698 => x"ff78f0c3",
  1699 => x"787148d4",
  1700 => x"c848d0ff",
  1701 => x"e0c078e1",
  1702 => x"0e4f2678",
  1703 => x"0e5c5b5e",
  1704 => x"f0c24c71",
  1705 => x"c6fc49e2",
  1706 => x"c04a7087",
  1707 => x"c204aab7",
  1708 => x"f0c387e2",
  1709 => x"87c905aa",
  1710 => x"48e0edc1",
  1711 => x"c3c278c1",
  1712 => x"aae0c387",
  1713 => x"c187c905",
  1714 => x"c148e4ed",
  1715 => x"87f4c178",
  1716 => x"bfe4edc1",
  1717 => x"c287c602",
  1718 => x"c24ba2c0",
  1719 => x"744b7287",
  1720 => x"87d1059c",
  1721 => x"bfe0edc1",
  1722 => x"e4edc11e",
  1723 => x"49721ebf",
  1724 => x"c887f9fd",
  1725 => x"e0edc186",
  1726 => x"e0c002bf",
  1727 => x"c4497387",
  1728 => x"c19129b7",
  1729 => x"7381c0ef",
  1730 => x"c29acf4a",
  1731 => x"7248c192",
  1732 => x"ff4a7030",
  1733 => x"694872ba",
  1734 => x"db797098",
  1735 => x"c4497387",
  1736 => x"c19129b7",
  1737 => x"7381c0ef",
  1738 => x"c29acf4a",
  1739 => x"7248c392",
  1740 => x"484a7030",
  1741 => x"7970b069",
  1742 => x"48e4edc1",
  1743 => x"edc178c0",
  1744 => x"78c048e0",
  1745 => x"49e2f0c2",
  1746 => x"7087e4f9",
  1747 => x"aab7c04a",
  1748 => x"87defd03",
  1749 => x"87c248c0",
  1750 => x"4c264d26",
  1751 => x"4f264b26",
  1752 => x"00000000",
  1753 => x"00000000",
  1754 => x"494a711e",
  1755 => x"2687ecfc",
  1756 => x"4ac01e4f",
  1757 => x"91c44972",
  1758 => x"81c0efc1",
  1759 => x"82c179c0",
  1760 => x"04aab7d0",
  1761 => x"4f2687ee",
  1762 => x"5c5b5e0e",
  1763 => x"4d710e5d",
  1764 => x"7587ccf8",
  1765 => x"2ab7c44a",
  1766 => x"c0efc192",
  1767 => x"cf4c7582",
  1768 => x"6a94c29c",
  1769 => x"2b744b49",
  1770 => x"48c29bc3",
  1771 => x"4c703074",
  1772 => x"4874bcff",
  1773 => x"7a709871",
  1774 => x"7387dcf7",
  1775 => x"87d8fe48",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"48d0ff1e",
  1793 => x"7178e1c8",
  1794 => x"08d4ff48",
  1795 => x"1e4f2678",
  1796 => x"c848d0ff",
  1797 => x"487178e1",
  1798 => x"7808d4ff",
  1799 => x"ff4866c4",
  1800 => x"267808d4",
  1801 => x"4a711e4f",
  1802 => x"1e4966c4",
  1803 => x"deff4972",
  1804 => x"48d0ff87",
  1805 => x"2678e0c0",
  1806 => x"731e4f26",
  1807 => x"c84b711e",
  1808 => x"731e4966",
  1809 => x"a2e0c14a",
  1810 => x"87d9ff49",
  1811 => x"2687c426",
  1812 => x"264c264d",
  1813 => x"1e4f264b",
  1814 => x"c34ad4ff",
  1815 => x"d0ff7aff",
  1816 => x"78e1c048",
  1817 => x"f0c27ade",
  1818 => x"497abfec",
  1819 => x"7028c848",
  1820 => x"d048717a",
  1821 => x"717a7028",
  1822 => x"7028d848",
  1823 => x"f0f0c27a",
  1824 => x"48497abf",
  1825 => x"7a7028c8",
  1826 => x"28d04871",
  1827 => x"48717a70",
  1828 => x"7a7028d8",
  1829 => x"c048d0ff",
  1830 => x"4f2678e0",
  1831 => x"711e731e",
  1832 => x"ecf0c24a",
  1833 => x"2b724bbf",
  1834 => x"04aae0c0",
  1835 => x"497287ce",
  1836 => x"c289e0c0",
  1837 => x"4bbff0f0",
  1838 => x"87cf2b71",
  1839 => x"7249e0c0",
  1840 => x"f0f0c289",
  1841 => x"307148bf",
  1842 => x"c8b34970",
  1843 => x"48739b66",
  1844 => x"4d2687c4",
  1845 => x"4b264c26",
  1846 => x"5e0e4f26",
  1847 => x"0e5d5c5b",
  1848 => x"4b7186ec",
  1849 => x"bfecf0c2",
  1850 => x"2c734c7e",
  1851 => x"04abe0c0",
  1852 => x"c487e0c0",
  1853 => x"78c048a6",
  1854 => x"e0c04973",
  1855 => x"c04a7189",
  1856 => x"724866e4",
  1857 => x"58a6cc30",
  1858 => x"bff0f0c2",
  1859 => x"2c714c4d",
  1860 => x"7387e4c0",
  1861 => x"66e4c049",
  1862 => x"c8307148",
  1863 => x"e0c058a6",
  1864 => x"c0897349",
  1865 => x"714866e4",
  1866 => x"58a6cc28",
  1867 => x"bff0f0c2",
  1868 => x"3071484d",
  1869 => x"c0b44970",
  1870 => x"c19c66e4",
  1871 => x"66e8c084",
  1872 => x"87c204ac",
  1873 => x"e0c04cc0",
  1874 => x"87d304ab",
  1875 => x"c048a6cc",
  1876 => x"c0497378",
  1877 => x"487489e0",
  1878 => x"a6d43071",
  1879 => x"7387d558",
  1880 => x"71487449",
  1881 => x"58a6d030",
  1882 => x"7349e0c0",
  1883 => x"71487489",
  1884 => x"58a6d428",
  1885 => x"ff4a66c4",
  1886 => x"c89a6eba",
  1887 => x"b9ff4966",
  1888 => x"48729975",
  1889 => x"c2b066cc",
  1890 => x"7158f0f0",
  1891 => x"b066d048",
  1892 => x"58f4f0c2",
  1893 => x"ec87c0fb",
  1894 => x"87f6fc8e",
  1895 => x"48d0ff1e",
  1896 => x"7178c9c8",
  1897 => x"08d4ff48",
  1898 => x"1e4f2678",
  1899 => x"eb494a71",
  1900 => x"48d0ff87",
  1901 => x"4f2678c8",
  1902 => x"711e731e",
  1903 => x"c0f1c24b",
  1904 => x"87c302bf",
  1905 => x"ff87ebc2",
  1906 => x"c9c848d0",
  1907 => x"c0497378",
  1908 => x"d4ffb1e0",
  1909 => x"c2787148",
  1910 => x"c048f4f0",
  1911 => x"0266c878",
  1912 => x"ffc387c5",
  1913 => x"c087c249",
  1914 => x"fcf0c249",
  1915 => x"0266cc59",
  1916 => x"d5c587c6",
  1917 => x"87c44ad5",
  1918 => x"4affffcf",
  1919 => x"5ac0f1c2",
  1920 => x"48c0f1c2",
  1921 => x"87c478c1",
  1922 => x"4c264d26",
  1923 => x"4f264b26",
  1924 => x"5c5b5e0e",
  1925 => x"4a710e5d",
  1926 => x"bffcf0c2",
  1927 => x"029a724c",
  1928 => x"c84987cb",
  1929 => x"eef6c191",
  1930 => x"c483714b",
  1931 => x"eefac187",
  1932 => x"134dc04b",
  1933 => x"c2997449",
  1934 => x"b9bff8f0",
  1935 => x"7148d4ff",
  1936 => x"2cb7c178",
  1937 => x"adb7c885",
  1938 => x"c287e804",
  1939 => x"48bff4f0",
  1940 => x"f0c280c8",
  1941 => x"effe58f8",
  1942 => x"1e731e87",
  1943 => x"4a134b71",
  1944 => x"87cb029a",
  1945 => x"e7fe4972",
  1946 => x"9a4a1387",
  1947 => x"fe87f505",
  1948 => x"c21e87da",
  1949 => x"49bff4f0",
  1950 => x"48f4f0c2",
  1951 => x"c478a1c1",
  1952 => x"03a9b7c0",
  1953 => x"d4ff87db",
  1954 => x"f8f0c248",
  1955 => x"f0c278bf",
  1956 => x"c249bff4",
  1957 => x"c148f4f0",
  1958 => x"c0c478a1",
  1959 => x"e504a9b7",
  1960 => x"48d0ff87",
  1961 => x"f1c278c8",
  1962 => x"78c048c0",
  1963 => x"00004f26",
  1964 => x"00000000",
  1965 => x"00000000",
  1966 => x"005f5f00",
  1967 => x"03000000",
  1968 => x"03030003",
  1969 => x"7f140000",
  1970 => x"7f7f147f",
  1971 => x"24000014",
  1972 => x"3a6b6b2e",
  1973 => x"6a4c0012",
  1974 => x"566c1836",
  1975 => x"7e300032",
  1976 => x"3a77594f",
  1977 => x"00004068",
  1978 => x"00030704",
  1979 => x"00000000",
  1980 => x"41633e1c",
  1981 => x"00000000",
  1982 => x"1c3e6341",
  1983 => x"2a080000",
  1984 => x"3e1c1c3e",
  1985 => x"0800082a",
  1986 => x"083e3e08",
  1987 => x"00000008",
  1988 => x"0060e080",
  1989 => x"08000000",
  1990 => x"08080808",
  1991 => x"00000008",
  1992 => x"00606000",
  1993 => x"60400000",
  1994 => x"060c1830",
  1995 => x"3e000103",
  1996 => x"7f4d597f",
  1997 => x"0400003e",
  1998 => x"007f7f06",
  1999 => x"42000000",
  2000 => x"4f597163",
  2001 => x"22000046",
  2002 => x"7f494963",
  2003 => x"1c180036",
  2004 => x"7f7f1316",
  2005 => x"27000010",
  2006 => x"7d454567",
  2007 => x"3c000039",
  2008 => x"79494b7e",
  2009 => x"01000030",
  2010 => x"0f797101",
  2011 => x"36000007",
  2012 => x"7f49497f",
  2013 => x"06000036",
  2014 => x"3f69494f",
  2015 => x"0000001e",
  2016 => x"00666600",
  2017 => x"00000000",
  2018 => x"0066e680",
  2019 => x"08000000",
  2020 => x"22141408",
  2021 => x"14000022",
  2022 => x"14141414",
  2023 => x"22000014",
  2024 => x"08141422",
  2025 => x"02000008",
  2026 => x"0f595103",
  2027 => x"7f3e0006",
  2028 => x"1f555d41",
  2029 => x"7e00001e",
  2030 => x"7f09097f",
  2031 => x"7f00007e",
  2032 => x"7f49497f",
  2033 => x"1c000036",
  2034 => x"4141633e",
  2035 => x"7f000041",
  2036 => x"3e63417f",
  2037 => x"7f00001c",
  2038 => x"4149497f",
  2039 => x"7f000041",
  2040 => x"0109097f",
  2041 => x"3e000001",
  2042 => x"7b49417f",
  2043 => x"7f00007a",
  2044 => x"7f08087f",
  2045 => x"0000007f",
  2046 => x"417f7f41",
  2047 => x"20000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
