library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"7f61417f",
     1 => x"0000407e",
     2 => x"19097f7f",
     3 => x"0000667f",
     4 => x"594d6f26",
     5 => x"0000327b",
     6 => x"7f7f0101",
     7 => x"00000101",
     8 => x"40407f3f",
     9 => x"00003f7f",
    10 => x"70703f0f",
    11 => x"7f000f3f",
    12 => x"3018307f",
    13 => x"41007f7f",
    14 => x"1c1c3663",
    15 => x"01416336",
    16 => x"7c7c0603",
    17 => x"61010306",
    18 => x"474d5971",
    19 => x"00004143",
    20 => x"417f7f00",
    21 => x"01000041",
    22 => x"180c0603",
    23 => x"00406030",
    24 => x"7f414100",
    25 => x"0800007f",
    26 => x"0603060c",
    27 => x"8000080c",
    28 => x"80808080",
    29 => x"00008080",
    30 => x"07030000",
    31 => x"00000004",
    32 => x"54547420",
    33 => x"0000787c",
    34 => x"44447f7f",
    35 => x"0000387c",
    36 => x"44447c38",
    37 => x"00000044",
    38 => x"44447c38",
    39 => x"00007f7f",
    40 => x"54547c38",
    41 => x"0000185c",
    42 => x"057f7e04",
    43 => x"00000005",
    44 => x"a4a4bc18",
    45 => x"00007cfc",
    46 => x"04047f7f",
    47 => x"0000787c",
    48 => x"7d3d0000",
    49 => x"00000040",
    50 => x"fd808080",
    51 => x"0000007d",
    52 => x"38107f7f",
    53 => x"0000446c",
    54 => x"7f3f0000",
    55 => x"7c000040",
    56 => x"0c180c7c",
    57 => x"0000787c",
    58 => x"04047c7c",
    59 => x"0000787c",
    60 => x"44447c38",
    61 => x"0000387c",
    62 => x"2424fcfc",
    63 => x"0000183c",
    64 => x"24243c18",
    65 => x"0000fcfc",
    66 => x"04047c7c",
    67 => x"0000080c",
    68 => x"54545c48",
    69 => x"00002074",
    70 => x"447f3f04",
    71 => x"00000044",
    72 => x"40407c3c",
    73 => x"00007c7c",
    74 => x"60603c1c",
    75 => x"3c001c3c",
    76 => x"6030607c",
    77 => x"44003c7c",
    78 => x"3810386c",
    79 => x"0000446c",
    80 => x"60e0bc1c",
    81 => x"00001c3c",
    82 => x"5c746444",
    83 => x"0000444c",
    84 => x"773e0808",
    85 => x"00004141",
    86 => x"7f7f0000",
    87 => x"00000000",
    88 => x"3e774141",
    89 => x"02000808",
    90 => x"02030101",
    91 => x"7f000102",
    92 => x"7f7f7f7f",
    93 => x"08007f7f",
    94 => x"3e1c1c08",
    95 => x"7f7f7f3e",
    96 => x"1c3e3e7f",
    97 => x"0008081c",
    98 => x"7c7c1810",
    99 => x"00001018",
   100 => x"7c7c3010",
   101 => x"10001030",
   102 => x"78606030",
   103 => x"4200061e",
   104 => x"3c183c66",
   105 => x"78004266",
   106 => x"c6c26a38",
   107 => x"6000386c",
   108 => x"00600000",
   109 => x"0e006000",
   110 => x"5d5c5b5e",
   111 => x"4c711e0e",
   112 => x"bfc1f1c2",
   113 => x"c04bc04d",
   114 => x"02ab741e",
   115 => x"a6c487c7",
   116 => x"c578c048",
   117 => x"48a6c487",
   118 => x"66c478c1",
   119 => x"ee49731e",
   120 => x"86c887df",
   121 => x"ef49e0c0",
   122 => x"a5c487ef",
   123 => x"f0496a4a",
   124 => x"c6f187f0",
   125 => x"c185cb87",
   126 => x"abb7c883",
   127 => x"87c7ff04",
   128 => x"264d2626",
   129 => x"264b264c",
   130 => x"4a711e4f",
   131 => x"5ac5f1c2",
   132 => x"48c5f1c2",
   133 => x"fe4978c7",
   134 => x"4f2687dd",
   135 => x"711e731e",
   136 => x"aab7c04a",
   137 => x"c287d303",
   138 => x"05bff6d5",
   139 => x"4bc187c4",
   140 => x"4bc087c2",
   141 => x"5bfad5c2",
   142 => x"d5c287c4",
   143 => x"d5c25afa",
   144 => x"c14abff6",
   145 => x"a2c0c19a",
   146 => x"87e8ec49",
   147 => x"d5c248fc",
   148 => x"fe78bff6",
   149 => x"711e87ef",
   150 => x"1e66c44a",
   151 => x"e2e64972",
   152 => x"4f262687",
   153 => x"f6d5c21e",
   154 => x"c4e349bf",
   155 => x"f9f0c287",
   156 => x"78bfe848",
   157 => x"48f5f0c2",
   158 => x"c278bfec",
   159 => x"4abff9f0",
   160 => x"99ffc349",
   161 => x"722ab7c8",
   162 => x"c2b07148",
   163 => x"2658c1f1",
   164 => x"5b5e0e4f",
   165 => x"710e5d5c",
   166 => x"87c8ff4b",
   167 => x"48f4f0c2",
   168 => x"497350c0",
   169 => x"7087eae2",
   170 => x"9cc24c49",
   171 => x"cb49eecb",
   172 => x"497087cc",
   173 => x"f4f0c24d",
   174 => x"c105bf97",
   175 => x"66d087e2",
   176 => x"fdf0c249",
   177 => x"d60599bf",
   178 => x"4966d487",
   179 => x"bff5f0c2",
   180 => x"87cb0599",
   181 => x"f8e14973",
   182 => x"02987087",
   183 => x"c187c1c1",
   184 => x"87c0fe4c",
   185 => x"e1ca4975",
   186 => x"02987087",
   187 => x"f0c287c6",
   188 => x"50c148f4",
   189 => x"97f4f0c2",
   190 => x"e3c005bf",
   191 => x"fdf0c287",
   192 => x"66d049bf",
   193 => x"d6ff0599",
   194 => x"f5f0c287",
   195 => x"66d449bf",
   196 => x"caff0599",
   197 => x"e0497387",
   198 => x"987087f7",
   199 => x"87fffe05",
   200 => x"dcfb4874",
   201 => x"5b5e0e87",
   202 => x"f40e5d5c",
   203 => x"4c4dc086",
   204 => x"c47ebfec",
   205 => x"f1c248a6",
   206 => x"c178bfc1",
   207 => x"c71ec01e",
   208 => x"87cdfd49",
   209 => x"987086c8",
   210 => x"ff87ce02",
   211 => x"87ccfb49",
   212 => x"ff49dac1",
   213 => x"c187fadf",
   214 => x"f4f0c24d",
   215 => x"c302bf97",
   216 => x"87c4d087",
   217 => x"bff9f0c2",
   218 => x"f6d5c24b",
   219 => x"ebc005bf",
   220 => x"49fdc387",
   221 => x"87d9dfff",
   222 => x"ff49fac3",
   223 => x"7387d2df",
   224 => x"99ffc349",
   225 => x"49c01e71",
   226 => x"7387cbfb",
   227 => x"29b7c849",
   228 => x"49c11e71",
   229 => x"c887fffa",
   230 => x"87c0c686",
   231 => x"bffdf0c2",
   232 => x"dd029b4b",
   233 => x"f2d5c287",
   234 => x"ddc749bf",
   235 => x"05987087",
   236 => x"4bc087c4",
   237 => x"e0c287d2",
   238 => x"87c2c749",
   239 => x"58f6d5c2",
   240 => x"d5c287c6",
   241 => x"78c048f2",
   242 => x"99c24973",
   243 => x"c387ce05",
   244 => x"ddff49eb",
   245 => x"497087fb",
   246 => x"c20299c2",
   247 => x"734cfb87",
   248 => x"0599c149",
   249 => x"f4c387ce",
   250 => x"e4ddff49",
   251 => x"c2497087",
   252 => x"87c20299",
   253 => x"49734cfa",
   254 => x"ce0599c8",
   255 => x"49f5c387",
   256 => x"87cdddff",
   257 => x"99c24970",
   258 => x"c287d502",
   259 => x"02bfc5f1",
   260 => x"c14887ca",
   261 => x"c9f1c288",
   262 => x"87c2c058",
   263 => x"4dc14cff",
   264 => x"99c44973",
   265 => x"c387ce05",
   266 => x"dcff49f2",
   267 => x"497087e3",
   268 => x"dc0299c2",
   269 => x"c5f1c287",
   270 => x"c7487ebf",
   271 => x"c003a8b7",
   272 => x"486e87cb",
   273 => x"f1c280c1",
   274 => x"c2c058c9",
   275 => x"c14cfe87",
   276 => x"49fdc34d",
   277 => x"87f9dbff",
   278 => x"99c24970",
   279 => x"c287d502",
   280 => x"02bfc5f1",
   281 => x"c287c9c0",
   282 => x"c048c5f1",
   283 => x"87c2c078",
   284 => x"4dc14cfd",
   285 => x"ff49fac3",
   286 => x"7087d6db",
   287 => x"0299c249",
   288 => x"c287d9c0",
   289 => x"48bfc5f1",
   290 => x"03a8b7c7",
   291 => x"c287c9c0",
   292 => x"c748c5f1",
   293 => x"87c2c078",
   294 => x"4dc14cfc",
   295 => x"03acb7c0",
   296 => x"c487d1c0",
   297 => x"d8c14a66",
   298 => x"c0026a82",
   299 => x"4b6a87c6",
   300 => x"0f734974",
   301 => x"f0c31ec0",
   302 => x"49dac11e",
   303 => x"c887d2f7",
   304 => x"02987086",
   305 => x"c887e2c0",
   306 => x"f1c248a6",
   307 => x"c878bfc5",
   308 => x"91cb4966",
   309 => x"714866c4",
   310 => x"6e7e7080",
   311 => x"c8c002bf",
   312 => x"4bbf6e87",
   313 => x"734966c8",
   314 => x"029d750f",
   315 => x"c287c8c0",
   316 => x"49bfc5f1",
   317 => x"c287c0f3",
   318 => x"02bffad5",
   319 => x"4987ddc0",
   320 => x"7087c7c2",
   321 => x"d3c00298",
   322 => x"c5f1c287",
   323 => x"e6f249bf",
   324 => x"f449c087",
   325 => x"d5c287c6",
   326 => x"78c048fa",
   327 => x"e0f38ef4",
   328 => x"5b5e0e87",
   329 => x"1e0e5d5c",
   330 => x"f1c24c71",
   331 => x"c149bfc1",
   332 => x"c14da1cd",
   333 => x"7e6981d1",
   334 => x"cf029c74",
   335 => x"4ba5c487",
   336 => x"f1c27b74",
   337 => x"f249bfc1",
   338 => x"7b6e87ff",
   339 => x"c4059c74",
   340 => x"c24bc087",
   341 => x"734bc187",
   342 => x"87c0f349",
   343 => x"c70266d4",
   344 => x"87da4987",
   345 => x"87c24a70",
   346 => x"d5c24ac0",
   347 => x"f2265afe",
   348 => x"000087cf",
   349 => x"00000000",
   350 => x"00000000",
   351 => x"711e0000",
   352 => x"bfc8ff4a",
   353 => x"48a17249",
   354 => x"ff1e4f26",
   355 => x"fe89bfc8",
   356 => x"c0c0c0c0",
   357 => x"c401a9c0",
   358 => x"c24ac087",
   359 => x"724ac187",
   360 => x"0e4f2648",
   361 => x"5d5c5b5e",
   362 => x"ff4b710e",
   363 => x"66d04cd4",
   364 => x"d678c048",
   365 => x"d0d8ff49",
   366 => x"7cffc387",
   367 => x"ffc3496c",
   368 => x"494d7199",
   369 => x"c199f0c3",
   370 => x"cb05a9e0",
   371 => x"7cffc387",
   372 => x"98c3486c",
   373 => x"780866d0",
   374 => x"6c7cffc3",
   375 => x"31c8494a",
   376 => x"6c7cffc3",
   377 => x"72b2714a",
   378 => x"c331c849",
   379 => x"4a6c7cff",
   380 => x"4972b271",
   381 => x"ffc331c8",
   382 => x"714a6c7c",
   383 => x"48d0ffb2",
   384 => x"7378e0c0",
   385 => x"87c2029b",
   386 => x"48757b72",
   387 => x"4c264d26",
   388 => x"4f264b26",
   389 => x"0e4f261e",
   390 => x"0e5c5b5e",
   391 => x"1e7686f8",
   392 => x"fd49a6c8",
   393 => x"86c487fd",
   394 => x"486e4b70",
   395 => x"c203a8c2",
   396 => x"4a7387f0",
   397 => x"c19af0c3",
   398 => x"c702aad0",
   399 => x"aae0c187",
   400 => x"87dec205",
   401 => x"99c84973",
   402 => x"ff87c302",
   403 => x"4c7387c6",
   404 => x"acc29cc3",
   405 => x"87c2c105",
   406 => x"c94966c4",
   407 => x"c41e7131",
   408 => x"92d44a66",
   409 => x"49c9f1c2",
   410 => x"cdfe8172",
   411 => x"49d887f2",
   412 => x"87d5d5ff",
   413 => x"c21ec0c8",
   414 => x"fd49e2df",
   415 => x"ff87ede9",
   416 => x"e0c048d0",
   417 => x"e2dfc278",
   418 => x"4a66cc1e",
   419 => x"f1c292d4",
   420 => x"817249c9",
   421 => x"87f9cbfe",
   422 => x"acc186cc",
   423 => x"87c2c105",
   424 => x"c94966c4",
   425 => x"c41e7131",
   426 => x"92d44a66",
   427 => x"49c9f1c2",
   428 => x"ccfe8172",
   429 => x"dfc287ea",
   430 => x"66c81ee2",
   431 => x"c292d44a",
   432 => x"7249c9f1",
   433 => x"f9c9fe81",
   434 => x"ff49d787",
   435 => x"c887fad3",
   436 => x"dfc21ec0",
   437 => x"e7fd49e2",
   438 => x"86cc87eb",
   439 => x"c048d0ff",
   440 => x"8ef878e0",
   441 => x"0e87e7fc",
   442 => x"5d5c5b5e",
   443 => x"4d711e0e",
   444 => x"d44cd4ff",
   445 => x"c3487e66",
   446 => x"c506a8b7",
   447 => x"c148c087",
   448 => x"497587e2",
   449 => x"87fedafe",
   450 => x"66c41e75",
   451 => x"c293d44b",
   452 => x"7383c9f1",
   453 => x"d4c5fe49",
   454 => x"6b83c887",
   455 => x"48d0ff4b",
   456 => x"dd78e1c8",
   457 => x"c349737c",
   458 => x"7c7199ff",
   459 => x"b7c84973",
   460 => x"99ffc329",
   461 => x"49737c71",
   462 => x"c329b7d0",
   463 => x"7c7199ff",
   464 => x"b7d84973",
   465 => x"c07c7129",
   466 => x"7c7c7c7c",
   467 => x"7c7c7c7c",
   468 => x"7c7c7c7c",
   469 => x"c478e0c0",
   470 => x"49dc1e66",
   471 => x"87ced2ff",
   472 => x"487386c8",
   473 => x"87e4fa26",
   474 => x"f6dec21e",
   475 => x"b9c149bf",
   476 => x"59fadec2",
   477 => x"c348d4ff",
   478 => x"d0ff78ff",
   479 => x"78e1c848",
   480 => x"c148d4ff",
   481 => x"7131c478",
   482 => x"48d0ff78",
   483 => x"2678e0c0",
   484 => x"dec21e4f",
   485 => x"ecc21eea",
   486 => x"c3fe49d8",
   487 => x"86c487cf",
   488 => x"c3029870",
   489 => x"87c0ff87",
   490 => x"35314f26",
   491 => x"205a484b",
   492 => x"46432020",
   493 => x"00000047",
   494 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
