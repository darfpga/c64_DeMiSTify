
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"7f",x"19",x"09",x"7f"),
     1 => (x"26",x"00",x"00",x"66"),
     2 => (x"7b",x"59",x"4d",x"6f"),
     3 => (x"01",x"00",x"00",x"32"),
     4 => (x"01",x"7f",x"7f",x"01"),
     5 => (x"3f",x"00",x"00",x"01"),
     6 => (x"7f",x"40",x"40",x"7f"),
     7 => (x"0f",x"00",x"00",x"3f"),
     8 => (x"3f",x"70",x"70",x"3f"),
     9 => (x"7f",x"7f",x"00",x"0f"),
    10 => (x"7f",x"30",x"18",x"30"),
    11 => (x"63",x"41",x"00",x"7f"),
    12 => (x"36",x"1c",x"1c",x"36"),
    13 => (x"03",x"01",x"41",x"63"),
    14 => (x"06",x"7c",x"7c",x"06"),
    15 => (x"71",x"61",x"01",x"03"),
    16 => (x"43",x"47",x"4d",x"59"),
    17 => (x"00",x"00",x"00",x"41"),
    18 => (x"41",x"41",x"7f",x"7f"),
    19 => (x"03",x"01",x"00",x"00"),
    20 => (x"30",x"18",x"0c",x"06"),
    21 => (x"00",x"00",x"40",x"60"),
    22 => (x"7f",x"7f",x"41",x"41"),
    23 => (x"0c",x"08",x"00",x"00"),
    24 => (x"0c",x"06",x"03",x"06"),
    25 => (x"80",x"80",x"00",x"08"),
    26 => (x"80",x"80",x"80",x"80"),
    27 => (x"00",x"00",x"00",x"80"),
    28 => (x"04",x"07",x"03",x"00"),
    29 => (x"20",x"00",x"00",x"00"),
    30 => (x"7c",x"54",x"54",x"74"),
    31 => (x"7f",x"00",x"00",x"78"),
    32 => (x"7c",x"44",x"44",x"7f"),
    33 => (x"38",x"00",x"00",x"38"),
    34 => (x"44",x"44",x"44",x"7c"),
    35 => (x"38",x"00",x"00",x"00"),
    36 => (x"7f",x"44",x"44",x"7c"),
    37 => (x"38",x"00",x"00",x"7f"),
    38 => (x"5c",x"54",x"54",x"7c"),
    39 => (x"04",x"00",x"00",x"18"),
    40 => (x"05",x"05",x"7f",x"7e"),
    41 => (x"18",x"00",x"00",x"00"),
    42 => (x"fc",x"a4",x"a4",x"bc"),
    43 => (x"7f",x"00",x"00",x"7c"),
    44 => (x"7c",x"04",x"04",x"7f"),
    45 => (x"00",x"00",x"00",x"78"),
    46 => (x"40",x"7d",x"3d",x"00"),
    47 => (x"80",x"00",x"00",x"00"),
    48 => (x"7d",x"fd",x"80",x"80"),
    49 => (x"7f",x"00",x"00",x"00"),
    50 => (x"6c",x"38",x"10",x"7f"),
    51 => (x"00",x"00",x"00",x"44"),
    52 => (x"40",x"7f",x"3f",x"00"),
    53 => (x"7c",x"7c",x"00",x"00"),
    54 => (x"7c",x"0c",x"18",x"0c"),
    55 => (x"7c",x"00",x"00",x"78"),
    56 => (x"7c",x"04",x"04",x"7c"),
    57 => (x"38",x"00",x"00",x"78"),
    58 => (x"7c",x"44",x"44",x"7c"),
    59 => (x"fc",x"00",x"00",x"38"),
    60 => (x"3c",x"24",x"24",x"fc"),
    61 => (x"18",x"00",x"00",x"18"),
    62 => (x"fc",x"24",x"24",x"3c"),
    63 => (x"7c",x"00",x"00",x"fc"),
    64 => (x"0c",x"04",x"04",x"7c"),
    65 => (x"48",x"00",x"00",x"08"),
    66 => (x"74",x"54",x"54",x"5c"),
    67 => (x"04",x"00",x"00",x"20"),
    68 => (x"44",x"44",x"7f",x"3f"),
    69 => (x"3c",x"00",x"00",x"00"),
    70 => (x"7c",x"40",x"40",x"7c"),
    71 => (x"1c",x"00",x"00",x"7c"),
    72 => (x"3c",x"60",x"60",x"3c"),
    73 => (x"7c",x"3c",x"00",x"1c"),
    74 => (x"7c",x"60",x"30",x"60"),
    75 => (x"6c",x"44",x"00",x"3c"),
    76 => (x"6c",x"38",x"10",x"38"),
    77 => (x"1c",x"00",x"00",x"44"),
    78 => (x"3c",x"60",x"e0",x"bc"),
    79 => (x"44",x"00",x"00",x"1c"),
    80 => (x"4c",x"5c",x"74",x"64"),
    81 => (x"08",x"00",x"00",x"44"),
    82 => (x"41",x"77",x"3e",x"08"),
    83 => (x"00",x"00",x"00",x"41"),
    84 => (x"00",x"7f",x"7f",x"00"),
    85 => (x"41",x"00",x"00",x"00"),
    86 => (x"08",x"3e",x"77",x"41"),
    87 => (x"01",x"02",x"00",x"08"),
    88 => (x"02",x"02",x"03",x"01"),
    89 => (x"7f",x"7f",x"00",x"01"),
    90 => (x"7f",x"7f",x"7f",x"7f"),
    91 => (x"08",x"08",x"00",x"7f"),
    92 => (x"3e",x"3e",x"1c",x"1c"),
    93 => (x"7f",x"7f",x"7f",x"7f"),
    94 => (x"1c",x"1c",x"3e",x"3e"),
    95 => (x"10",x"00",x"08",x"08"),
    96 => (x"18",x"7c",x"7c",x"18"),
    97 => (x"10",x"00",x"00",x"10"),
    98 => (x"30",x"7c",x"7c",x"30"),
    99 => (x"30",x"10",x"00",x"10"),
   100 => (x"1e",x"78",x"60",x"60"),
   101 => (x"66",x"42",x"00",x"06"),
   102 => (x"66",x"3c",x"18",x"3c"),
   103 => (x"38",x"78",x"00",x"42"),
   104 => (x"6c",x"c6",x"c2",x"6a"),
   105 => (x"00",x"60",x"00",x"38"),
   106 => (x"00",x"00",x"60",x"00"),
   107 => (x"5e",x"0e",x"00",x"60"),
   108 => (x"0e",x"5d",x"5c",x"5b"),
   109 => (x"c2",x"4c",x"71",x"1e"),
   110 => (x"4d",x"bf",x"d1",x"f0"),
   111 => (x"1e",x"c0",x"4b",x"c0"),
   112 => (x"c7",x"02",x"ab",x"74"),
   113 => (x"48",x"a6",x"c4",x"87"),
   114 => (x"87",x"c5",x"78",x"c0"),
   115 => (x"c1",x"48",x"a6",x"c4"),
   116 => (x"1e",x"66",x"c4",x"78"),
   117 => (x"df",x"ee",x"49",x"73"),
   118 => (x"c0",x"86",x"c8",x"87"),
   119 => (x"ef",x"ef",x"49",x"e0"),
   120 => (x"4a",x"a5",x"c4",x"87"),
   121 => (x"f0",x"f0",x"49",x"6a"),
   122 => (x"87",x"c6",x"f1",x"87"),
   123 => (x"83",x"c1",x"85",x"cb"),
   124 => (x"04",x"ab",x"b7",x"c8"),
   125 => (x"26",x"87",x"c7",x"ff"),
   126 => (x"4c",x"26",x"4d",x"26"),
   127 => (x"4f",x"26",x"4b",x"26"),
   128 => (x"c2",x"4a",x"71",x"1e"),
   129 => (x"c2",x"5a",x"d5",x"f0"),
   130 => (x"c7",x"48",x"d5",x"f0"),
   131 => (x"dd",x"fe",x"49",x"78"),
   132 => (x"1e",x"4f",x"26",x"87"),
   133 => (x"4a",x"71",x"1e",x"73"),
   134 => (x"03",x"aa",x"b7",x"c0"),
   135 => (x"d5",x"c2",x"87",x"d3"),
   136 => (x"c4",x"05",x"bf",x"ed"),
   137 => (x"c2",x"4b",x"c1",x"87"),
   138 => (x"c2",x"4b",x"c0",x"87"),
   139 => (x"c4",x"5b",x"f1",x"d5"),
   140 => (x"f1",x"d5",x"c2",x"87"),
   141 => (x"ed",x"d5",x"c2",x"5a"),
   142 => (x"9a",x"c1",x"4a",x"bf"),
   143 => (x"49",x"a2",x"c0",x"c1"),
   144 => (x"fc",x"87",x"e8",x"ec"),
   145 => (x"ed",x"d5",x"c2",x"48"),
   146 => (x"ef",x"fe",x"78",x"bf"),
   147 => (x"4a",x"71",x"1e",x"87"),
   148 => (x"72",x"1e",x"66",x"c4"),
   149 => (x"87",x"e2",x"e6",x"49"),
   150 => (x"1e",x"4f",x"26",x"26"),
   151 => (x"bf",x"ed",x"d5",x"c2"),
   152 => (x"87",x"c4",x"e3",x"49"),
   153 => (x"48",x"c9",x"f0",x"c2"),
   154 => (x"c2",x"78",x"bf",x"e8"),
   155 => (x"ec",x"48",x"c5",x"f0"),
   156 => (x"f0",x"c2",x"78",x"bf"),
   157 => (x"49",x"4a",x"bf",x"c9"),
   158 => (x"c8",x"99",x"ff",x"c3"),
   159 => (x"48",x"72",x"2a",x"b7"),
   160 => (x"f0",x"c2",x"b0",x"71"),
   161 => (x"4f",x"26",x"58",x"d1"),
   162 => (x"5c",x"5b",x"5e",x"0e"),
   163 => (x"4b",x"71",x"0e",x"5d"),
   164 => (x"c2",x"87",x"c8",x"ff"),
   165 => (x"c0",x"48",x"c4",x"f0"),
   166 => (x"e2",x"49",x"73",x"50"),
   167 => (x"49",x"70",x"87",x"ea"),
   168 => (x"cb",x"9c",x"c2",x"4c"),
   169 => (x"cc",x"cb",x"49",x"ee"),
   170 => (x"4d",x"49",x"70",x"87"),
   171 => (x"97",x"c4",x"f0",x"c2"),
   172 => (x"e2",x"c1",x"05",x"bf"),
   173 => (x"49",x"66",x"d0",x"87"),
   174 => (x"bf",x"cd",x"f0",x"c2"),
   175 => (x"87",x"d6",x"05",x"99"),
   176 => (x"c2",x"49",x"66",x"d4"),
   177 => (x"99",x"bf",x"c5",x"f0"),
   178 => (x"73",x"87",x"cb",x"05"),
   179 => (x"87",x"f8",x"e1",x"49"),
   180 => (x"c1",x"02",x"98",x"70"),
   181 => (x"4c",x"c1",x"87",x"c1"),
   182 => (x"75",x"87",x"c0",x"fe"),
   183 => (x"87",x"e1",x"ca",x"49"),
   184 => (x"c6",x"02",x"98",x"70"),
   185 => (x"c4",x"f0",x"c2",x"87"),
   186 => (x"c2",x"50",x"c1",x"48"),
   187 => (x"bf",x"97",x"c4",x"f0"),
   188 => (x"87",x"e3",x"c0",x"05"),
   189 => (x"bf",x"cd",x"f0",x"c2"),
   190 => (x"99",x"66",x"d0",x"49"),
   191 => (x"87",x"d6",x"ff",x"05"),
   192 => (x"bf",x"c5",x"f0",x"c2"),
   193 => (x"99",x"66",x"d4",x"49"),
   194 => (x"87",x"ca",x"ff",x"05"),
   195 => (x"f7",x"e0",x"49",x"73"),
   196 => (x"05",x"98",x"70",x"87"),
   197 => (x"74",x"87",x"ff",x"fe"),
   198 => (x"87",x"dc",x"fb",x"48"),
   199 => (x"5c",x"5b",x"5e",x"0e"),
   200 => (x"86",x"f4",x"0e",x"5d"),
   201 => (x"ec",x"4c",x"4d",x"c0"),
   202 => (x"a6",x"c4",x"7e",x"bf"),
   203 => (x"d1",x"f0",x"c2",x"48"),
   204 => (x"1e",x"c1",x"78",x"bf"),
   205 => (x"49",x"c7",x"1e",x"c0"),
   206 => (x"c8",x"87",x"cd",x"fd"),
   207 => (x"02",x"98",x"70",x"86"),
   208 => (x"49",x"ff",x"87",x"ce"),
   209 => (x"c1",x"87",x"cc",x"fb"),
   210 => (x"df",x"ff",x"49",x"da"),
   211 => (x"4d",x"c1",x"87",x"fa"),
   212 => (x"97",x"c4",x"f0",x"c2"),
   213 => (x"87",x"c3",x"02",x"bf"),
   214 => (x"c2",x"87",x"c4",x"d0"),
   215 => (x"4b",x"bf",x"c9",x"f0"),
   216 => (x"bf",x"ed",x"d5",x"c2"),
   217 => (x"87",x"eb",x"c0",x"05"),
   218 => (x"ff",x"49",x"fd",x"c3"),
   219 => (x"c3",x"87",x"d9",x"df"),
   220 => (x"df",x"ff",x"49",x"fa"),
   221 => (x"49",x"73",x"87",x"d2"),
   222 => (x"71",x"99",x"ff",x"c3"),
   223 => (x"fb",x"49",x"c0",x"1e"),
   224 => (x"49",x"73",x"87",x"cb"),
   225 => (x"71",x"29",x"b7",x"c8"),
   226 => (x"fa",x"49",x"c1",x"1e"),
   227 => (x"86",x"c8",x"87",x"ff"),
   228 => (x"c2",x"87",x"c0",x"c6"),
   229 => (x"4b",x"bf",x"cd",x"f0"),
   230 => (x"87",x"dd",x"02",x"9b"),
   231 => (x"bf",x"e9",x"d5",x"c2"),
   232 => (x"87",x"dd",x"c7",x"49"),
   233 => (x"c4",x"05",x"98",x"70"),
   234 => (x"d2",x"4b",x"c0",x"87"),
   235 => (x"49",x"e0",x"c2",x"87"),
   236 => (x"c2",x"87",x"c2",x"c7"),
   237 => (x"c6",x"58",x"ed",x"d5"),
   238 => (x"e9",x"d5",x"c2",x"87"),
   239 => (x"73",x"78",x"c0",x"48"),
   240 => (x"05",x"99",x"c2",x"49"),
   241 => (x"eb",x"c3",x"87",x"ce"),
   242 => (x"fb",x"dd",x"ff",x"49"),
   243 => (x"c2",x"49",x"70",x"87"),
   244 => (x"87",x"c2",x"02",x"99"),
   245 => (x"49",x"73",x"4c",x"fb"),
   246 => (x"ce",x"05",x"99",x"c1"),
   247 => (x"49",x"f4",x"c3",x"87"),
   248 => (x"87",x"e4",x"dd",x"ff"),
   249 => (x"99",x"c2",x"49",x"70"),
   250 => (x"fa",x"87",x"c2",x"02"),
   251 => (x"c8",x"49",x"73",x"4c"),
   252 => (x"87",x"ce",x"05",x"99"),
   253 => (x"ff",x"49",x"f5",x"c3"),
   254 => (x"70",x"87",x"cd",x"dd"),
   255 => (x"02",x"99",x"c2",x"49"),
   256 => (x"f0",x"c2",x"87",x"d5"),
   257 => (x"ca",x"02",x"bf",x"d5"),
   258 => (x"88",x"c1",x"48",x"87"),
   259 => (x"58",x"d9",x"f0",x"c2"),
   260 => (x"ff",x"87",x"c2",x"c0"),
   261 => (x"73",x"4d",x"c1",x"4c"),
   262 => (x"05",x"99",x"c4",x"49"),
   263 => (x"f2",x"c3",x"87",x"ce"),
   264 => (x"e3",x"dc",x"ff",x"49"),
   265 => (x"c2",x"49",x"70",x"87"),
   266 => (x"87",x"dc",x"02",x"99"),
   267 => (x"bf",x"d5",x"f0",x"c2"),
   268 => (x"b7",x"c7",x"48",x"7e"),
   269 => (x"cb",x"c0",x"03",x"a8"),
   270 => (x"c1",x"48",x"6e",x"87"),
   271 => (x"d9",x"f0",x"c2",x"80"),
   272 => (x"87",x"c2",x"c0",x"58"),
   273 => (x"4d",x"c1",x"4c",x"fe"),
   274 => (x"ff",x"49",x"fd",x"c3"),
   275 => (x"70",x"87",x"f9",x"db"),
   276 => (x"02",x"99",x"c2",x"49"),
   277 => (x"f0",x"c2",x"87",x"d5"),
   278 => (x"c0",x"02",x"bf",x"d5"),
   279 => (x"f0",x"c2",x"87",x"c9"),
   280 => (x"78",x"c0",x"48",x"d5"),
   281 => (x"fd",x"87",x"c2",x"c0"),
   282 => (x"c3",x"4d",x"c1",x"4c"),
   283 => (x"db",x"ff",x"49",x"fa"),
   284 => (x"49",x"70",x"87",x"d6"),
   285 => (x"c0",x"02",x"99",x"c2"),
   286 => (x"f0",x"c2",x"87",x"d9"),
   287 => (x"c7",x"48",x"bf",x"d5"),
   288 => (x"c0",x"03",x"a8",x"b7"),
   289 => (x"f0",x"c2",x"87",x"c9"),
   290 => (x"78",x"c7",x"48",x"d5"),
   291 => (x"fc",x"87",x"c2",x"c0"),
   292 => (x"c0",x"4d",x"c1",x"4c"),
   293 => (x"c0",x"03",x"ac",x"b7"),
   294 => (x"66",x"c4",x"87",x"d1"),
   295 => (x"82",x"d8",x"c1",x"4a"),
   296 => (x"c6",x"c0",x"02",x"6a"),
   297 => (x"74",x"4b",x"6a",x"87"),
   298 => (x"c0",x"0f",x"73",x"49"),
   299 => (x"1e",x"f0",x"c3",x"1e"),
   300 => (x"f7",x"49",x"da",x"c1"),
   301 => (x"86",x"c8",x"87",x"d2"),
   302 => (x"c0",x"02",x"98",x"70"),
   303 => (x"a6",x"c8",x"87",x"e2"),
   304 => (x"d5",x"f0",x"c2",x"48"),
   305 => (x"66",x"c8",x"78",x"bf"),
   306 => (x"c4",x"91",x"cb",x"49"),
   307 => (x"80",x"71",x"48",x"66"),
   308 => (x"bf",x"6e",x"7e",x"70"),
   309 => (x"87",x"c8",x"c0",x"02"),
   310 => (x"c8",x"4b",x"bf",x"6e"),
   311 => (x"0f",x"73",x"49",x"66"),
   312 => (x"c0",x"02",x"9d",x"75"),
   313 => (x"f0",x"c2",x"87",x"c8"),
   314 => (x"f3",x"49",x"bf",x"d5"),
   315 => (x"d5",x"c2",x"87",x"c0"),
   316 => (x"c0",x"02",x"bf",x"f1"),
   317 => (x"c2",x"49",x"87",x"dd"),
   318 => (x"98",x"70",x"87",x"c7"),
   319 => (x"87",x"d3",x"c0",x"02"),
   320 => (x"bf",x"d5",x"f0",x"c2"),
   321 => (x"87",x"e6",x"f2",x"49"),
   322 => (x"c6",x"f4",x"49",x"c0"),
   323 => (x"f1",x"d5",x"c2",x"87"),
   324 => (x"f4",x"78",x"c0",x"48"),
   325 => (x"87",x"e0",x"f3",x"8e"),
   326 => (x"5c",x"5b",x"5e",x"0e"),
   327 => (x"71",x"1e",x"0e",x"5d"),
   328 => (x"d1",x"f0",x"c2",x"4c"),
   329 => (x"cd",x"c1",x"49",x"bf"),
   330 => (x"d1",x"c1",x"4d",x"a1"),
   331 => (x"74",x"7e",x"69",x"81"),
   332 => (x"87",x"cf",x"02",x"9c"),
   333 => (x"74",x"4b",x"a5",x"c4"),
   334 => (x"d1",x"f0",x"c2",x"7b"),
   335 => (x"ff",x"f2",x"49",x"bf"),
   336 => (x"74",x"7b",x"6e",x"87"),
   337 => (x"87",x"c4",x"05",x"9c"),
   338 => (x"87",x"c2",x"4b",x"c0"),
   339 => (x"49",x"73",x"4b",x"c1"),
   340 => (x"d4",x"87",x"c0",x"f3"),
   341 => (x"87",x"c7",x"02",x"66"),
   342 => (x"70",x"87",x"da",x"49"),
   343 => (x"c0",x"87",x"c2",x"4a"),
   344 => (x"f5",x"d5",x"c2",x"4a"),
   345 => (x"cf",x"f2",x"26",x"5a"),
   346 => (x"00",x"00",x"00",x"87"),
   347 => (x"00",x"00",x"00",x"00"),
   348 => (x"00",x"00",x"00",x"00"),
   349 => (x"4a",x"71",x"1e",x"00"),
   350 => (x"49",x"bf",x"c8",x"ff"),
   351 => (x"26",x"48",x"a1",x"72"),
   352 => (x"c8",x"ff",x"1e",x"4f"),
   353 => (x"c0",x"fe",x"89",x"bf"),
   354 => (x"c0",x"c0",x"c0",x"c0"),
   355 => (x"87",x"c4",x"01",x"a9"),
   356 => (x"87",x"c2",x"4a",x"c0"),
   357 => (x"48",x"72",x"4a",x"c1"),
   358 => (x"5e",x"0e",x"4f",x"26"),
   359 => (x"0e",x"5d",x"5c",x"5b"),
   360 => (x"d4",x"ff",x"4b",x"71"),
   361 => (x"48",x"66",x"d0",x"4c"),
   362 => (x"49",x"d6",x"78",x"c0"),
   363 => (x"87",x"d0",x"d8",x"ff"),
   364 => (x"6c",x"7c",x"ff",x"c3"),
   365 => (x"99",x"ff",x"c3",x"49"),
   366 => (x"c3",x"49",x"4d",x"71"),
   367 => (x"e0",x"c1",x"99",x"f0"),
   368 => (x"87",x"cb",x"05",x"a9"),
   369 => (x"6c",x"7c",x"ff",x"c3"),
   370 => (x"d0",x"98",x"c3",x"48"),
   371 => (x"c3",x"78",x"08",x"66"),
   372 => (x"4a",x"6c",x"7c",x"ff"),
   373 => (x"c3",x"31",x"c8",x"49"),
   374 => (x"4a",x"6c",x"7c",x"ff"),
   375 => (x"49",x"72",x"b2",x"71"),
   376 => (x"ff",x"c3",x"31",x"c8"),
   377 => (x"71",x"4a",x"6c",x"7c"),
   378 => (x"c8",x"49",x"72",x"b2"),
   379 => (x"7c",x"ff",x"c3",x"31"),
   380 => (x"b2",x"71",x"4a",x"6c"),
   381 => (x"c0",x"48",x"d0",x"ff"),
   382 => (x"9b",x"73",x"78",x"e0"),
   383 => (x"72",x"87",x"c2",x"02"),
   384 => (x"26",x"48",x"75",x"7b"),
   385 => (x"26",x"4c",x"26",x"4d"),
   386 => (x"1e",x"4f",x"26",x"4b"),
   387 => (x"5e",x"0e",x"4f",x"26"),
   388 => (x"f8",x"0e",x"5c",x"5b"),
   389 => (x"c8",x"1e",x"76",x"86"),
   390 => (x"fd",x"fd",x"49",x"a6"),
   391 => (x"70",x"86",x"c4",x"87"),
   392 => (x"c2",x"48",x"6e",x"4b"),
   393 => (x"f0",x"c2",x"03",x"a8"),
   394 => (x"c3",x"4a",x"73",x"87"),
   395 => (x"d0",x"c1",x"9a",x"f0"),
   396 => (x"87",x"c7",x"02",x"aa"),
   397 => (x"05",x"aa",x"e0",x"c1"),
   398 => (x"73",x"87",x"de",x"c2"),
   399 => (x"02",x"99",x"c8",x"49"),
   400 => (x"c6",x"ff",x"87",x"c3"),
   401 => (x"c3",x"4c",x"73",x"87"),
   402 => (x"05",x"ac",x"c2",x"9c"),
   403 => (x"c4",x"87",x"c2",x"c1"),
   404 => (x"31",x"c9",x"49",x"66"),
   405 => (x"66",x"c4",x"1e",x"71"),
   406 => (x"c2",x"92",x"d4",x"4a"),
   407 => (x"72",x"49",x"d9",x"f0"),
   408 => (x"fb",x"cd",x"fe",x"81"),
   409 => (x"ff",x"49",x"d8",x"87"),
   410 => (x"c8",x"87",x"d5",x"d5"),
   411 => (x"de",x"c2",x"1e",x"c0"),
   412 => (x"e9",x"fd",x"49",x"f2"),
   413 => (x"d0",x"ff",x"87",x"f6"),
   414 => (x"78",x"e0",x"c0",x"48"),
   415 => (x"1e",x"f2",x"de",x"c2"),
   416 => (x"d4",x"4a",x"66",x"cc"),
   417 => (x"d9",x"f0",x"c2",x"92"),
   418 => (x"fe",x"81",x"72",x"49"),
   419 => (x"cc",x"87",x"c2",x"cc"),
   420 => (x"05",x"ac",x"c1",x"86"),
   421 => (x"c4",x"87",x"c2",x"c1"),
   422 => (x"31",x"c9",x"49",x"66"),
   423 => (x"66",x"c4",x"1e",x"71"),
   424 => (x"c2",x"92",x"d4",x"4a"),
   425 => (x"72",x"49",x"d9",x"f0"),
   426 => (x"f3",x"cc",x"fe",x"81"),
   427 => (x"f2",x"de",x"c2",x"87"),
   428 => (x"4a",x"66",x"c8",x"1e"),
   429 => (x"f0",x"c2",x"92",x"d4"),
   430 => (x"81",x"72",x"49",x"d9"),
   431 => (x"87",x"c2",x"ca",x"fe"),
   432 => (x"d3",x"ff",x"49",x"d7"),
   433 => (x"c0",x"c8",x"87",x"fa"),
   434 => (x"f2",x"de",x"c2",x"1e"),
   435 => (x"f4",x"e7",x"fd",x"49"),
   436 => (x"ff",x"86",x"cc",x"87"),
   437 => (x"e0",x"c0",x"48",x"d0"),
   438 => (x"fc",x"8e",x"f8",x"78"),
   439 => (x"5e",x"0e",x"87",x"e7"),
   440 => (x"0e",x"5d",x"5c",x"5b"),
   441 => (x"ff",x"4d",x"71",x"1e"),
   442 => (x"66",x"d4",x"4c",x"d4"),
   443 => (x"b7",x"c3",x"48",x"7e"),
   444 => (x"87",x"c5",x"06",x"a8"),
   445 => (x"e2",x"c1",x"48",x"c0"),
   446 => (x"fe",x"49",x"75",x"87"),
   447 => (x"75",x"87",x"c7",x"db"),
   448 => (x"4b",x"66",x"c4",x"1e"),
   449 => (x"f0",x"c2",x"93",x"d4"),
   450 => (x"49",x"73",x"83",x"d9"),
   451 => (x"87",x"fe",x"c3",x"fe"),
   452 => (x"4b",x"6b",x"83",x"c8"),
   453 => (x"c8",x"48",x"d0",x"ff"),
   454 => (x"7c",x"dd",x"78",x"e1"),
   455 => (x"ff",x"c3",x"49",x"73"),
   456 => (x"73",x"7c",x"71",x"99"),
   457 => (x"29",x"b7",x"c8",x"49"),
   458 => (x"71",x"99",x"ff",x"c3"),
   459 => (x"d0",x"49",x"73",x"7c"),
   460 => (x"ff",x"c3",x"29",x"b7"),
   461 => (x"73",x"7c",x"71",x"99"),
   462 => (x"29",x"b7",x"d8",x"49"),
   463 => (x"7c",x"c0",x"7c",x"71"),
   464 => (x"7c",x"7c",x"7c",x"7c"),
   465 => (x"7c",x"7c",x"7c",x"7c"),
   466 => (x"c0",x"7c",x"7c",x"7c"),
   467 => (x"66",x"c4",x"78",x"e0"),
   468 => (x"ff",x"49",x"dc",x"1e"),
   469 => (x"c8",x"87",x"ce",x"d2"),
   470 => (x"26",x"48",x"73",x"86"),
   471 => (x"1e",x"87",x"e4",x"fa"),
   472 => (x"bf",x"c8",x"de",x"c2"),
   473 => (x"c2",x"b9",x"c1",x"49"),
   474 => (x"ff",x"59",x"cc",x"de"),
   475 => (x"ff",x"c3",x"48",x"d4"),
   476 => (x"48",x"d0",x"ff",x"78"),
   477 => (x"ff",x"78",x"e1",x"c0"),
   478 => (x"78",x"c1",x"48",x"d4"),
   479 => (x"78",x"71",x"31",x"c4"),
   480 => (x"c0",x"48",x"d0",x"ff"),
   481 => (x"4f",x"26",x"78",x"e0"),
   482 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

