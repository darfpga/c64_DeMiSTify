library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"ccf2c287",
    12 => x"86c0c84e",
    13 => x"49ccf2c2",
    14 => x"48d4dfc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087dfe2",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"c44a711e",
    47 => x"c1484966",
    48 => x"58a6c888",
    49 => x"d4029971",
    50 => x"ff481287",
    51 => x"c47808d4",
    52 => x"c1484966",
    53 => x"58a6c888",
    54 => x"ec059971",
    55 => x"1e4f2687",
    56 => x"66c44a71",
    57 => x"88c14849",
    58 => x"7158a6c8",
    59 => x"87d60299",
    60 => x"c348d4ff",
    61 => x"526878ff",
    62 => x"484966c4",
    63 => x"a6c888c1",
    64 => x"05997158",
    65 => x"4f2687ea",
    66 => x"ff1e731e",
    67 => x"ffc34bd4",
    68 => x"c34a6b7b",
    69 => x"496b7bff",
    70 => x"b17232c8",
    71 => x"6b7bffc3",
    72 => x"7131c84a",
    73 => x"7bffc3b2",
    74 => x"32c8496b",
    75 => x"4871b172",
    76 => x"4d2687c4",
    77 => x"4b264c26",
    78 => x"5e0e4f26",
    79 => x"0e5d5c5b",
    80 => x"d4ff4a71",
    81 => x"c349724c",
    82 => x"7c7199ff",
    83 => x"bfd4dfc2",
    84 => x"d087c805",
    85 => x"30c94866",
    86 => x"d058a6d4",
    87 => x"29d84966",
    88 => x"7199ffc3",
    89 => x"4966d07c",
    90 => x"ffc329d0",
    91 => x"d07c7199",
    92 => x"29c84966",
    93 => x"7199ffc3",
    94 => x"4966d07c",
    95 => x"7199ffc3",
    96 => x"d049727c",
    97 => x"99ffc329",
    98 => x"4b6c7c71",
    99 => x"4dfff0c9",
   100 => x"05abffc3",
   101 => x"ffc387d0",
   102 => x"c14b6c7c",
   103 => x"87c6028d",
   104 => x"02abffc3",
   105 => x"487387f0",
   106 => x"1e87c7fe",
   107 => x"d4ff49c0",
   108 => x"78ffc348",
   109 => x"c8c381c1",
   110 => x"f104a9b7",
   111 => x"1e4f2687",
   112 => x"87e71e73",
   113 => x"4bdff8c4",
   114 => x"ffc01ec0",
   115 => x"49f7c1f0",
   116 => x"c487e7fd",
   117 => x"05a8c186",
   118 => x"ff87eac0",
   119 => x"ffc348d4",
   120 => x"c0c0c178",
   121 => x"1ec0c0c0",
   122 => x"c1f0e1c0",
   123 => x"c9fd49e9",
   124 => x"7086c487",
   125 => x"87ca0598",
   126 => x"c348d4ff",
   127 => x"48c178ff",
   128 => x"e6fe87cb",
   129 => x"058bc187",
   130 => x"c087fdfe",
   131 => x"87e6fc48",
   132 => x"ff1e731e",
   133 => x"ffc348d4",
   134 => x"c04bd378",
   135 => x"f0ffc01e",
   136 => x"fc49c1c1",
   137 => x"86c487d4",
   138 => x"ca059870",
   139 => x"48d4ff87",
   140 => x"c178ffc3",
   141 => x"fd87cb48",
   142 => x"8bc187f1",
   143 => x"87dbff05",
   144 => x"f1fb48c0",
   145 => x"5b5e0e87",
   146 => x"d4ff0e5c",
   147 => x"87dbfd4c",
   148 => x"c01eeac6",
   149 => x"c8c1f0e1",
   150 => x"87defb49",
   151 => x"a8c186c4",
   152 => x"fe87c802",
   153 => x"48c087ea",
   154 => x"fa87e2c1",
   155 => x"497087da",
   156 => x"99ffffcf",
   157 => x"02a9eac6",
   158 => x"d3fe87c8",
   159 => x"c148c087",
   160 => x"ffc387cb",
   161 => x"4bf1c07c",
   162 => x"7087f4fc",
   163 => x"ebc00298",
   164 => x"c01ec087",
   165 => x"fac1f0ff",
   166 => x"87defa49",
   167 => x"987086c4",
   168 => x"c387d905",
   169 => x"496c7cff",
   170 => x"7c7cffc3",
   171 => x"c0c17c7c",
   172 => x"87c40299",
   173 => x"87d548c1",
   174 => x"87d148c0",
   175 => x"c405abc2",
   176 => x"c848c087",
   177 => x"058bc187",
   178 => x"c087fdfe",
   179 => x"87e4f948",
   180 => x"c21e731e",
   181 => x"c148d4df",
   182 => x"ff4bc778",
   183 => x"78c248d0",
   184 => x"ff87c8fb",
   185 => x"78c348d0",
   186 => x"e5c01ec0",
   187 => x"49c0c1d0",
   188 => x"c487c7f9",
   189 => x"05a8c186",
   190 => x"c24b87c1",
   191 => x"87c505ab",
   192 => x"f9c048c0",
   193 => x"058bc187",
   194 => x"fc87d0ff",
   195 => x"dfc287f7",
   196 => x"987058d8",
   197 => x"c187cd05",
   198 => x"f0ffc01e",
   199 => x"f849d0c1",
   200 => x"86c487d8",
   201 => x"c348d4ff",
   202 => x"dec478ff",
   203 => x"dcdfc287",
   204 => x"48d0ff58",
   205 => x"d4ff78c2",
   206 => x"78ffc348",
   207 => x"f5f748c1",
   208 => x"5b5e0e87",
   209 => x"710e5d5c",
   210 => x"4dffc34a",
   211 => x"754cd4ff",
   212 => x"48d0ff7c",
   213 => x"7578c3c4",
   214 => x"c01e727c",
   215 => x"d8c1f0ff",
   216 => x"87d6f749",
   217 => x"987086c4",
   218 => x"c187c502",
   219 => x"87f0c048",
   220 => x"fec37c75",
   221 => x"1ec0c87c",
   222 => x"f44966d4",
   223 => x"86c487fa",
   224 => x"7c757c75",
   225 => x"dad87c75",
   226 => x"7c754be0",
   227 => x"0599496c",
   228 => x"8bc187c5",
   229 => x"7587f305",
   230 => x"48d0ff7c",
   231 => x"48c078c2",
   232 => x"0e87cff6",
   233 => x"5d5c5b5e",
   234 => x"c04b710e",
   235 => x"cdeec54c",
   236 => x"d4ff4adf",
   237 => x"78ffc348",
   238 => x"fec34968",
   239 => x"fdc005a9",
   240 => x"734d7087",
   241 => x"87cc029b",
   242 => x"731e66d0",
   243 => x"87cff449",
   244 => x"87d686c4",
   245 => x"c448d0ff",
   246 => x"ffc378d1",
   247 => x"4866d07d",
   248 => x"a6d488c1",
   249 => x"05987058",
   250 => x"d4ff87f0",
   251 => x"78ffc348",
   252 => x"059b7378",
   253 => x"d0ff87c5",
   254 => x"c178d048",
   255 => x"8ac14c4a",
   256 => x"87eefe05",
   257 => x"e9f44874",
   258 => x"1e731e87",
   259 => x"4bc04a71",
   260 => x"c348d4ff",
   261 => x"d0ff78ff",
   262 => x"78c3c448",
   263 => x"c348d4ff",
   264 => x"1e7278ff",
   265 => x"c1f0ffc0",
   266 => x"cdf449d1",
   267 => x"7086c487",
   268 => x"87d20598",
   269 => x"cc1ec0c8",
   270 => x"e6fd4966",
   271 => x"7086c487",
   272 => x"48d0ff4b",
   273 => x"487378c2",
   274 => x"0e87ebf3",
   275 => x"5d5c5b5e",
   276 => x"c01ec00e",
   277 => x"c9c1f0ff",
   278 => x"87def349",
   279 => x"dfc21ed2",
   280 => x"fefc49dc",
   281 => x"c086c887",
   282 => x"d284c14c",
   283 => x"f804acb7",
   284 => x"dcdfc287",
   285 => x"c349bf97",
   286 => x"c0c199c0",
   287 => x"e7c005a9",
   288 => x"e3dfc287",
   289 => x"d049bf97",
   290 => x"e4dfc231",
   291 => x"c84abf97",
   292 => x"c2b17232",
   293 => x"bf97e5df",
   294 => x"4c71b14a",
   295 => x"ffffffcf",
   296 => x"ca84c19c",
   297 => x"87e7c134",
   298 => x"97e5dfc2",
   299 => x"31c149bf",
   300 => x"dfc299c6",
   301 => x"4abf97e6",
   302 => x"722ab7c7",
   303 => x"e1dfc2b1",
   304 => x"4d4abf97",
   305 => x"dfc29dcf",
   306 => x"4abf97e2",
   307 => x"32ca9ac3",
   308 => x"97e3dfc2",
   309 => x"33c24bbf",
   310 => x"dfc2b273",
   311 => x"4bbf97e4",
   312 => x"c69bc0c3",
   313 => x"b2732bb7",
   314 => x"48c181c2",
   315 => x"49703071",
   316 => x"307548c1",
   317 => x"4c724d70",
   318 => x"947184c1",
   319 => x"adb7c0c8",
   320 => x"c187cc06",
   321 => x"c82db734",
   322 => x"01adb7c0",
   323 => x"7487f4ff",
   324 => x"87def048",
   325 => x"5c5b5e0e",
   326 => x"86f80e5d",
   327 => x"48c2e8c2",
   328 => x"dfc278c0",
   329 => x"49c01efa",
   330 => x"c487defb",
   331 => x"05987086",
   332 => x"48c087c5",
   333 => x"c087cec9",
   334 => x"c07ec14d",
   335 => x"49bff6f2",
   336 => x"4af0e0c2",
   337 => x"ec4bc871",
   338 => x"987087e0",
   339 => x"c087c205",
   340 => x"f2f2c07e",
   341 => x"e1c249bf",
   342 => x"c8714acc",
   343 => x"87caec4b",
   344 => x"c2059870",
   345 => x"6e7ec087",
   346 => x"87fdc002",
   347 => x"bfc0e7c2",
   348 => x"f8e7c24d",
   349 => x"487ebf9f",
   350 => x"a8ead6c5",
   351 => x"c287c705",
   352 => x"4dbfc0e7",
   353 => x"486e87ce",
   354 => x"a8d5e9ca",
   355 => x"c087c502",
   356 => x"87f1c748",
   357 => x"1efadfc2",
   358 => x"ecf94975",
   359 => x"7086c487",
   360 => x"87c50598",
   361 => x"dcc748c0",
   362 => x"f2f2c087",
   363 => x"e1c249bf",
   364 => x"c8714acc",
   365 => x"87f2ea4b",
   366 => x"c8059870",
   367 => x"c2e8c287",
   368 => x"da78c148",
   369 => x"f6f2c087",
   370 => x"e0c249bf",
   371 => x"c8714af0",
   372 => x"87d6ea4b",
   373 => x"c0029870",
   374 => x"48c087c5",
   375 => x"c287e6c6",
   376 => x"bf97f8e7",
   377 => x"a9d5c149",
   378 => x"87cdc005",
   379 => x"97f9e7c2",
   380 => x"eac249bf",
   381 => x"c5c002a9",
   382 => x"c648c087",
   383 => x"dfc287c7",
   384 => x"7ebf97fa",
   385 => x"a8e9c348",
   386 => x"87cec002",
   387 => x"ebc3486e",
   388 => x"c5c002a8",
   389 => x"c548c087",
   390 => x"e0c287eb",
   391 => x"49bf97c5",
   392 => x"ccc00599",
   393 => x"c6e0c287",
   394 => x"c249bf97",
   395 => x"c5c002a9",
   396 => x"c548c087",
   397 => x"e0c287cf",
   398 => x"48bf97c7",
   399 => x"58fee7c2",
   400 => x"c1484c70",
   401 => x"c2e8c288",
   402 => x"c8e0c258",
   403 => x"7549bf97",
   404 => x"c9e0c281",
   405 => x"c84abf97",
   406 => x"7ea17232",
   407 => x"48cfecc2",
   408 => x"e0c2786e",
   409 => x"48bf97ca",
   410 => x"c258a6c8",
   411 => x"02bfc2e8",
   412 => x"c087d4c2",
   413 => x"49bff2f2",
   414 => x"4acce1c2",
   415 => x"e74bc871",
   416 => x"987087e8",
   417 => x"87c5c002",
   418 => x"f8c348c0",
   419 => x"fae7c287",
   420 => x"ecc24cbf",
   421 => x"e0c25ce3",
   422 => x"49bf97df",
   423 => x"e0c231c8",
   424 => x"4abf97de",
   425 => x"e0c249a1",
   426 => x"4abf97e0",
   427 => x"a17232d0",
   428 => x"e1e0c249",
   429 => x"d84abf97",
   430 => x"49a17232",
   431 => x"c29166c4",
   432 => x"81bfcfec",
   433 => x"59d7ecc2",
   434 => x"97e7e0c2",
   435 => x"32c84abf",
   436 => x"97e6e0c2",
   437 => x"4aa24bbf",
   438 => x"97e8e0c2",
   439 => x"33d04bbf",
   440 => x"c24aa273",
   441 => x"bf97e9e0",
   442 => x"d89bcf4b",
   443 => x"4aa27333",
   444 => x"5adbecc2",
   445 => x"bfd7ecc2",
   446 => x"748ac24a",
   447 => x"dbecc292",
   448 => x"78a17248",
   449 => x"c287cac1",
   450 => x"bf97cce0",
   451 => x"c231c849",
   452 => x"bf97cbe0",
   453 => x"c249a14a",
   454 => x"c259cae8",
   455 => x"49bfc6e8",
   456 => x"ffc731c5",
   457 => x"c229c981",
   458 => x"c259e3ec",
   459 => x"bf97d1e0",
   460 => x"c232c84a",
   461 => x"bf97d0e0",
   462 => x"c44aa24b",
   463 => x"826e9266",
   464 => x"5adfecc2",
   465 => x"48d7ecc2",
   466 => x"ecc278c0",
   467 => x"a17248d3",
   468 => x"e3ecc278",
   469 => x"d7ecc248",
   470 => x"ecc278bf",
   471 => x"ecc248e7",
   472 => x"c278bfdb",
   473 => x"02bfc2e8",
   474 => x"7487c9c0",
   475 => x"7030c448",
   476 => x"87c9c07e",
   477 => x"bfdfecc2",
   478 => x"7030c448",
   479 => x"c6e8c27e",
   480 => x"c1786e48",
   481 => x"268ef848",
   482 => x"264c264d",
   483 => x"0e4f264b",
   484 => x"5d5c5b5e",
   485 => x"c24a710e",
   486 => x"02bfc2e8",
   487 => x"4b7287cb",
   488 => x"4c722bc7",
   489 => x"c99cffc1",
   490 => x"c84b7287",
   491 => x"c34c722b",
   492 => x"ecc29cff",
   493 => x"c083bfcf",
   494 => x"abbfeef2",
   495 => x"c087d902",
   496 => x"c25bf2f2",
   497 => x"731efadf",
   498 => x"87fdf049",
   499 => x"987086c4",
   500 => x"c087c505",
   501 => x"87e6c048",
   502 => x"bfc2e8c2",
   503 => x"7487d202",
   504 => x"c291c449",
   505 => x"6981fadf",
   506 => x"ffffcf4d",
   507 => x"cb9dffff",
   508 => x"c2497487",
   509 => x"fadfc291",
   510 => x"4d699f81",
   511 => x"c6fe4875",
   512 => x"5b5e0e87",
   513 => x"f80e5d5c",
   514 => x"9c4c7186",
   515 => x"c087c505",
   516 => x"87c1c348",
   517 => x"6e7ea4c8",
   518 => x"d878c048",
   519 => x"87c70266",
   520 => x"bf9766d8",
   521 => x"c087c505",
   522 => x"87e9c248",
   523 => x"49c11ec0",
   524 => x"c487e0ca",
   525 => x"9d4d7086",
   526 => x"87c2c102",
   527 => x"4acae8c2",
   528 => x"e04966d8",
   529 => x"987087c9",
   530 => x"87f2c002",
   531 => x"66d84a75",
   532 => x"e04bcb49",
   533 => x"987087ee",
   534 => x"87e2c002",
   535 => x"9d751ec0",
   536 => x"c887c702",
   537 => x"78c048a6",
   538 => x"a6c887c5",
   539 => x"c878c148",
   540 => x"dec94966",
   541 => x"7086c487",
   542 => x"fe059d4d",
   543 => x"9d7587fe",
   544 => x"87cfc102",
   545 => x"6e49a5dc",
   546 => x"da786948",
   547 => x"a6c449a5",
   548 => x"78a4c448",
   549 => x"c448699f",
   550 => x"c2780866",
   551 => x"02bfc2e8",
   552 => x"a5d487d2",
   553 => x"49699f49",
   554 => x"99ffffc0",
   555 => x"30d04871",
   556 => x"87c27e70",
   557 => x"496e7ec0",
   558 => x"bf66c448",
   559 => x"0866c480",
   560 => x"cc7cc078",
   561 => x"66c449a4",
   562 => x"a4d079bf",
   563 => x"c179c049",
   564 => x"c087c248",
   565 => x"fa8ef848",
   566 => x"5e0e87ed",
   567 => x"0e5d5c5b",
   568 => x"029c4c71",
   569 => x"c887cac1",
   570 => x"026949a4",
   571 => x"d087c2c1",
   572 => x"496c4a66",
   573 => x"5aa6d482",
   574 => x"b94d66d0",
   575 => x"bffee7c2",
   576 => x"72baff4a",
   577 => x"02997199",
   578 => x"c487e4c0",
   579 => x"496b4ba4",
   580 => x"7087fcf9",
   581 => x"fae7c27b",
   582 => x"816c49bf",
   583 => x"b9757c71",
   584 => x"bffee7c2",
   585 => x"72baff4a",
   586 => x"05997199",
   587 => x"7587dcff",
   588 => x"87d3f97c",
   589 => x"711e731e",
   590 => x"c7029b4b",
   591 => x"49a3c887",
   592 => x"87c50569",
   593 => x"f7c048c0",
   594 => x"d3ecc287",
   595 => x"a3c44abf",
   596 => x"c2496949",
   597 => x"fae7c289",
   598 => x"a27191bf",
   599 => x"fee7c24a",
   600 => x"996b49bf",
   601 => x"c04aa271",
   602 => x"c85af2f2",
   603 => x"49721e66",
   604 => x"c487d6ea",
   605 => x"05987086",
   606 => x"48c087c4",
   607 => x"48c187c2",
   608 => x"1e87c8f8",
   609 => x"4b711e73",
   610 => x"87c7029b",
   611 => x"6949a3c8",
   612 => x"c087c505",
   613 => x"87f7c048",
   614 => x"bfd3ecc2",
   615 => x"49a3c44a",
   616 => x"89c24969",
   617 => x"bffae7c2",
   618 => x"4aa27191",
   619 => x"bffee7c2",
   620 => x"71996b49",
   621 => x"f2c04aa2",
   622 => x"66c85af2",
   623 => x"e549721e",
   624 => x"86c487ff",
   625 => x"c4059870",
   626 => x"c248c087",
   627 => x"f648c187",
   628 => x"5e0e87f9",
   629 => x"1e0e5c5b",
   630 => x"66d04b71",
   631 => x"732cc94c",
   632 => x"d4c1029b",
   633 => x"49a3c887",
   634 => x"ccc10269",
   635 => x"fee7c287",
   636 => x"b9ff49bf",
   637 => x"7e994a6b",
   638 => x"d103ac71",
   639 => x"d07bc087",
   640 => x"79c049a3",
   641 => x"c44aa3cc",
   642 => x"796a49a3",
   643 => x"8c7287c2",
   644 => x"c0029c74",
   645 => x"1e4987e3",
   646 => x"fdfa4973",
   647 => x"d086c487",
   648 => x"ffc74966",
   649 => x"87cb0299",
   650 => x"1efadfc2",
   651 => x"c3fc4973",
   652 => x"d086c487",
   653 => x"66d049a3",
   654 => x"ccf52679",
   655 => x"1e731e87",
   656 => x"029b4b71",
   657 => x"c287e4c0",
   658 => x"735be7ec",
   659 => x"c28ac24a",
   660 => x"49bffae7",
   661 => x"d3ecc292",
   662 => x"807248bf",
   663 => x"58ebecc2",
   664 => x"30c44871",
   665 => x"58cae8c2",
   666 => x"c287edc0",
   667 => x"c248e3ec",
   668 => x"78bfd7ec",
   669 => x"48e7ecc2",
   670 => x"bfdbecc2",
   671 => x"c2e8c278",
   672 => x"87c902bf",
   673 => x"bffae7c2",
   674 => x"c731c449",
   675 => x"dfecc287",
   676 => x"31c449bf",
   677 => x"59cae8c2",
   678 => x"0e87f0f3",
   679 => x"0e5c5b5e",
   680 => x"4bc04a71",
   681 => x"c0029a72",
   682 => x"a2da87e1",
   683 => x"4b699f49",
   684 => x"bfc2e8c2",
   685 => x"d487cf02",
   686 => x"699f49a2",
   687 => x"ffc04c49",
   688 => x"34d09cff",
   689 => x"4cc087c2",
   690 => x"73b34974",
   691 => x"87edfd49",
   692 => x"0e87f6f2",
   693 => x"5d5c5b5e",
   694 => x"7186f40e",
   695 => x"727ec04a",
   696 => x"87d8029a",
   697 => x"48f6dfc2",
   698 => x"dfc278c0",
   699 => x"ecc248ee",
   700 => x"c278bfe7",
   701 => x"c248f2df",
   702 => x"78bfe3ec",
   703 => x"48d7e8c2",
   704 => x"e8c250c0",
   705 => x"c249bfc6",
   706 => x"4abff6df",
   707 => x"c403aa71",
   708 => x"497287c9",
   709 => x"c00599cf",
   710 => x"f2c087e9",
   711 => x"dfc248ee",
   712 => x"c278bfee",
   713 => x"c21efadf",
   714 => x"49bfeedf",
   715 => x"48eedfc2",
   716 => x"7178a1c1",
   717 => x"c487d2e3",
   718 => x"eaf2c086",
   719 => x"fadfc248",
   720 => x"c087cc78",
   721 => x"48bfeaf2",
   722 => x"c080e0c0",
   723 => x"c258eef2",
   724 => x"48bff6df",
   725 => x"dfc280c1",
   726 => x"aa2758fa",
   727 => x"bf00000c",
   728 => x"9d4dbf97",
   729 => x"87e3c202",
   730 => x"02ade5c3",
   731 => x"c087dcc2",
   732 => x"4bbfeaf2",
   733 => x"1149a3cb",
   734 => x"05accf4c",
   735 => x"7587d2c1",
   736 => x"c199df49",
   737 => x"c291cd89",
   738 => x"c181cae8",
   739 => x"51124aa3",
   740 => x"124aa3c3",
   741 => x"4aa3c551",
   742 => x"a3c75112",
   743 => x"c951124a",
   744 => x"51124aa3",
   745 => x"124aa3ce",
   746 => x"4aa3d051",
   747 => x"a3d25112",
   748 => x"d451124a",
   749 => x"51124aa3",
   750 => x"124aa3d6",
   751 => x"4aa3d851",
   752 => x"a3dc5112",
   753 => x"de51124a",
   754 => x"51124aa3",
   755 => x"fac07ec1",
   756 => x"c8497487",
   757 => x"ebc00599",
   758 => x"d0497487",
   759 => x"87d10599",
   760 => x"c00266dc",
   761 => x"497387cb",
   762 => x"700f66dc",
   763 => x"d3c00298",
   764 => x"c0056e87",
   765 => x"e8c287c6",
   766 => x"50c048ca",
   767 => x"bfeaf2c0",
   768 => x"87e1c248",
   769 => x"48d7e8c2",
   770 => x"c27e50c0",
   771 => x"49bfc6e8",
   772 => x"bff6dfc2",
   773 => x"04aa714a",
   774 => x"c287f7fb",
   775 => x"05bfe7ec",
   776 => x"c287c8c0",
   777 => x"02bfc2e8",
   778 => x"c287f8c1",
   779 => x"49bff2df",
   780 => x"7087dced",
   781 => x"f6dfc249",
   782 => x"48a6c459",
   783 => x"bff2dfc2",
   784 => x"c2e8c278",
   785 => x"d8c002bf",
   786 => x"4966c487",
   787 => x"ffffffcf",
   788 => x"02a999f8",
   789 => x"c087c5c0",
   790 => x"87e1c04c",
   791 => x"dcc04cc1",
   792 => x"4966c487",
   793 => x"99f8ffcf",
   794 => x"c8c002a9",
   795 => x"48a6c887",
   796 => x"c5c078c0",
   797 => x"48a6c887",
   798 => x"66c878c1",
   799 => x"059c744c",
   800 => x"c487e0c0",
   801 => x"89c24966",
   802 => x"bffae7c2",
   803 => x"ecc2914a",
   804 => x"c24abfd3",
   805 => x"7248eedf",
   806 => x"dfc278a1",
   807 => x"78c048f6",
   808 => x"c087dff9",
   809 => x"eb8ef448",
   810 => x"000087dd",
   811 => x"ffff0000",
   812 => x"0cbaffff",
   813 => x"0cc30000",
   814 => x"41460000",
   815 => x"20323354",
   816 => x"46002020",
   817 => x"36315441",
   818 => x"00202020",
   819 => x"48d4ff1e",
   820 => x"6878ffc3",
   821 => x"1e4f2648",
   822 => x"c348d4ff",
   823 => x"d0ff78ff",
   824 => x"78e1c048",
   825 => x"d448d4ff",
   826 => x"ebecc278",
   827 => x"bfd4ff48",
   828 => x"1e4f2650",
   829 => x"c048d0ff",
   830 => x"4f2678e0",
   831 => x"87ccff1e",
   832 => x"02994970",
   833 => x"fbc087c6",
   834 => x"87f105a9",
   835 => x"4f264871",
   836 => x"5c5b5e0e",
   837 => x"c04b710e",
   838 => x"87f0fe4c",
   839 => x"02994970",
   840 => x"c087f9c0",
   841 => x"c002a9ec",
   842 => x"fbc087f2",
   843 => x"ebc002a9",
   844 => x"b766cc87",
   845 => x"87c703ac",
   846 => x"c20266d0",
   847 => x"71537187",
   848 => x"87c20299",
   849 => x"c3fe84c1",
   850 => x"99497087",
   851 => x"c087cd02",
   852 => x"c702a9ec",
   853 => x"a9fbc087",
   854 => x"87d5ff05",
   855 => x"c30266d0",
   856 => x"7b97c087",
   857 => x"05a9ecc0",
   858 => x"4a7487c4",
   859 => x"4a7487c5",
   860 => x"728a0ac0",
   861 => x"2687c248",
   862 => x"264c264d",
   863 => x"1e4f264b",
   864 => x"7087c9fd",
   865 => x"f0c04a49",
   866 => x"87c904aa",
   867 => x"01aaf9c0",
   868 => x"f0c087c3",
   869 => x"aac1c18a",
   870 => x"c187c904",
   871 => x"c301aada",
   872 => x"8af7c087",
   873 => x"04aae1c1",
   874 => x"fac187c9",
   875 => x"87c301aa",
   876 => x"728afdc0",
   877 => x"0e4f2648",
   878 => x"0e5c5b5e",
   879 => x"d4ff4a71",
   880 => x"c049724c",
   881 => x"4b7087e9",
   882 => x"87c2029b",
   883 => x"d0ff8bc1",
   884 => x"c178c548",
   885 => x"49737cd5",
   886 => x"e4c131c6",
   887 => x"4abf97c0",
   888 => x"70b07148",
   889 => x"48d0ff7c",
   890 => x"487378c4",
   891 => x"0e87cafe",
   892 => x"5d5c5b5e",
   893 => x"7186f80e",
   894 => x"fb7ec04c",
   895 => x"4bc087d9",
   896 => x"97dcfac0",
   897 => x"a9c049bf",
   898 => x"fb87cf04",
   899 => x"83c187ee",
   900 => x"97dcfac0",
   901 => x"06ab49bf",
   902 => x"fac087f1",
   903 => x"02bf97dc",
   904 => x"e7fa87cf",
   905 => x"99497087",
   906 => x"c087c602",
   907 => x"f105a9ec",
   908 => x"fa4bc087",
   909 => x"4d7087d6",
   910 => x"c887d1fa",
   911 => x"cbfa58a6",
   912 => x"c14a7087",
   913 => x"49a4c883",
   914 => x"ad496997",
   915 => x"c087c702",
   916 => x"c005adff",
   917 => x"a4c987e7",
   918 => x"49699749",
   919 => x"02a966c4",
   920 => x"c04887c7",
   921 => x"d405a8ff",
   922 => x"49a4ca87",
   923 => x"aa496997",
   924 => x"c087c602",
   925 => x"c405aaff",
   926 => x"d07ec187",
   927 => x"adecc087",
   928 => x"c087c602",
   929 => x"c405adfb",
   930 => x"c14bc087",
   931 => x"fe026e7e",
   932 => x"def987e1",
   933 => x"f8487387",
   934 => x"87dbfb8e",
   935 => x"5b5e0e00",
   936 => x"f80e5d5c",
   937 => x"ff4d7186",
   938 => x"1e754bd4",
   939 => x"49f0ecc2",
   940 => x"c487cee5",
   941 => x"02987086",
   942 => x"c487d2c4",
   943 => x"e4c148a6",
   944 => x"7578bfc2",
   945 => x"87effb49",
   946 => x"c548d0ff",
   947 => x"7bd6c178",
   948 => x"a2754ac0",
   949 => x"c17b1149",
   950 => x"aab7cb82",
   951 => x"cc87f304",
   952 => x"7bffc34a",
   953 => x"e0c082c1",
   954 => x"f404aab7",
   955 => x"48d0ff87",
   956 => x"ffc378c4",
   957 => x"c178c57b",
   958 => x"7bc17bd3",
   959 => x"486678c4",
   960 => x"06a8b7c0",
   961 => x"c287f6c2",
   962 => x"4cbff8ec",
   963 => x"744866c4",
   964 => x"58a6c888",
   965 => x"c1029c74",
   966 => x"dfc287ff",
   967 => x"c0c87efa",
   968 => x"b7c08c4d",
   969 => x"87c603ac",
   970 => x"4da4c0c8",
   971 => x"c0c84cc0",
   972 => x"87dc05ad",
   973 => x"97ebecc2",
   974 => x"99d049bf",
   975 => x"c087d102",
   976 => x"f0ecc21e",
   977 => x"87ece749",
   978 => x"497086c4",
   979 => x"87eec04a",
   980 => x"1efadfc2",
   981 => x"49f0ecc2",
   982 => x"c487d9e7",
   983 => x"4a497086",
   984 => x"c848d0ff",
   985 => x"d4c178c5",
   986 => x"bf976e7b",
   987 => x"c1486e7b",
   988 => x"c17e7080",
   989 => x"f0ff058d",
   990 => x"48d0ff87",
   991 => x"9a7278c4",
   992 => x"c087c505",
   993 => x"87c7c148",
   994 => x"ecc21ec1",
   995 => x"c9e549f0",
   996 => x"7486c487",
   997 => x"c1fe059c",
   998 => x"4866c487",
   999 => x"06a8b7c0",
  1000 => x"ecc287d1",
  1001 => x"78c048f0",
  1002 => x"78c080d0",
  1003 => x"ecc280f4",
  1004 => x"c478bffc",
  1005 => x"b7c04866",
  1006 => x"cafd01a8",
  1007 => x"48d0ff87",
  1008 => x"d3c178c5",
  1009 => x"c47bc07b",
  1010 => x"c248c178",
  1011 => x"f848c087",
  1012 => x"264d268e",
  1013 => x"264b264c",
  1014 => x"5b5e0e4f",
  1015 => x"1e0e5d5c",
  1016 => x"4cc04b71",
  1017 => x"c004ab4d",
  1018 => x"f7c087e8",
  1019 => x"9d751eef",
  1020 => x"c087c402",
  1021 => x"c187c24a",
  1022 => x"eb49724a",
  1023 => x"86c487d5",
  1024 => x"84c17e70",
  1025 => x"87c2056e",
  1026 => x"85c14c73",
  1027 => x"ff06ac73",
  1028 => x"486e87d8",
  1029 => x"87f9fe26",
  1030 => x"5c5b5e0e",
  1031 => x"cc4b710e",
  1032 => x"87d80266",
  1033 => x"8cf0c04c",
  1034 => x"7487d802",
  1035 => x"028ac14a",
  1036 => x"028a87d1",
  1037 => x"028a87cd",
  1038 => x"87d987c9",
  1039 => x"dcf94973",
  1040 => x"7487d287",
  1041 => x"c149c01e",
  1042 => x"7487d9db",
  1043 => x"c149731e",
  1044 => x"c887d1db",
  1045 => x"87fbfd86",
  1046 => x"5c5b5e0e",
  1047 => x"711e0e5d",
  1048 => x"91de494c",
  1049 => x"4dd8edc2",
  1050 => x"6d978571",
  1051 => x"87dcc102",
  1052 => x"bfc4edc2",
  1053 => x"7282744a",
  1054 => x"87ddfd49",
  1055 => x"026e7e70",
  1056 => x"c287f2c0",
  1057 => x"6e4bcced",
  1058 => x"ff49cb4a",
  1059 => x"7487d9c0",
  1060 => x"c193cb4b",
  1061 => x"c483d4e4",
  1062 => x"d0c3c183",
  1063 => x"c149747b",
  1064 => x"7587d1c5",
  1065 => x"c1e4c17b",
  1066 => x"1e49bf97",
  1067 => x"49ccedc2",
  1068 => x"c487e5fd",
  1069 => x"c1497486",
  1070 => x"c087f9c4",
  1071 => x"d8c6c149",
  1072 => x"ececc287",
  1073 => x"c178c048",
  1074 => x"87d9dd49",
  1075 => x"87c1fc26",
  1076 => x"64616f4c",
  1077 => x"2e676e69",
  1078 => x"0e002e2e",
  1079 => x"0e5c5b5e",
  1080 => x"c24a4b71",
  1081 => x"82bfc4ed",
  1082 => x"ecfb4972",
  1083 => x"9c4c7087",
  1084 => x"4987c402",
  1085 => x"c287e4e6",
  1086 => x"c048c4ed",
  1087 => x"dc49c178",
  1088 => x"cefb87e3",
  1089 => x"5b5e0e87",
  1090 => x"f40e5d5c",
  1091 => x"fadfc286",
  1092 => x"c44cc04d",
  1093 => x"78c048a6",
  1094 => x"bfc4edc2",
  1095 => x"06a9c049",
  1096 => x"c287c1c1",
  1097 => x"9848fadf",
  1098 => x"87f8c002",
  1099 => x"1eeff7c0",
  1100 => x"c70266c8",
  1101 => x"48a6c487",
  1102 => x"87c578c0",
  1103 => x"c148a6c4",
  1104 => x"4966c478",
  1105 => x"c487cce6",
  1106 => x"c14d7086",
  1107 => x"4866c484",
  1108 => x"a6c880c1",
  1109 => x"c4edc258",
  1110 => x"03ac49bf",
  1111 => x"9d7587c6",
  1112 => x"87c8ff05",
  1113 => x"9d754cc0",
  1114 => x"87e0c302",
  1115 => x"1eeff7c0",
  1116 => x"c70266c8",
  1117 => x"48a6cc87",
  1118 => x"87c578c0",
  1119 => x"c148a6cc",
  1120 => x"4966cc78",
  1121 => x"c487cce5",
  1122 => x"6e7e7086",
  1123 => x"87e9c202",
  1124 => x"81cb496e",
  1125 => x"d0496997",
  1126 => x"d6c10299",
  1127 => x"dbc3c187",
  1128 => x"cb49744a",
  1129 => x"d4e4c191",
  1130 => x"c8797281",
  1131 => x"51ffc381",
  1132 => x"91de4974",
  1133 => x"4dd8edc2",
  1134 => x"c1c28571",
  1135 => x"a5c17d97",
  1136 => x"51e0c049",
  1137 => x"97cae8c2",
  1138 => x"87d202bf",
  1139 => x"a5c284c1",
  1140 => x"cae8c24b",
  1141 => x"fe49db4a",
  1142 => x"c187cdfb",
  1143 => x"a5cd87db",
  1144 => x"c151c049",
  1145 => x"4ba5c284",
  1146 => x"49cb4a6e",
  1147 => x"87f8fafe",
  1148 => x"c187c6c1",
  1149 => x"744ad8c1",
  1150 => x"c191cb49",
  1151 => x"7281d4e4",
  1152 => x"cae8c279",
  1153 => x"d802bf97",
  1154 => x"de497487",
  1155 => x"c284c191",
  1156 => x"714bd8ed",
  1157 => x"cae8c283",
  1158 => x"fe49dd4a",
  1159 => x"d887c9fa",
  1160 => x"de4b7487",
  1161 => x"d8edc293",
  1162 => x"49a3cb83",
  1163 => x"84c151c0",
  1164 => x"cb4a6e73",
  1165 => x"eff9fe49",
  1166 => x"4866c487",
  1167 => x"a6c880c1",
  1168 => x"03acc758",
  1169 => x"6e87c5c0",
  1170 => x"87e0fc05",
  1171 => x"8ef44874",
  1172 => x"1e87fef5",
  1173 => x"4b711e73",
  1174 => x"c191cb49",
  1175 => x"c881d4e4",
  1176 => x"e4c14aa1",
  1177 => x"501248c0",
  1178 => x"c04aa1c9",
  1179 => x"1248dcfa",
  1180 => x"c181ca50",
  1181 => x"1148c1e4",
  1182 => x"c1e4c150",
  1183 => x"1e49bf97",
  1184 => x"d3f649c0",
  1185 => x"ececc287",
  1186 => x"c178de48",
  1187 => x"87d5d649",
  1188 => x"87c1f526",
  1189 => x"494a711e",
  1190 => x"e4c191cb",
  1191 => x"81c881d4",
  1192 => x"ecc24811",
  1193 => x"edc258f0",
  1194 => x"78c048c4",
  1195 => x"f4d549c1",
  1196 => x"1e4f2687",
  1197 => x"fec049c0",
  1198 => x"4f2687df",
  1199 => x"0299711e",
  1200 => x"e5c187d2",
  1201 => x"50c048e9",
  1202 => x"cac180f7",
  1203 => x"e4c140d4",
  1204 => x"87ce78cd",
  1205 => x"48e5e5c1",
  1206 => x"78c6e4c1",
  1207 => x"cac180fc",
  1208 => x"4f2678f3",
  1209 => x"5c5b5e0e",
  1210 => x"4a4c710e",
  1211 => x"e4c192cb",
  1212 => x"a2c882d4",
  1213 => x"4ba2c949",
  1214 => x"1e4b6b97",
  1215 => x"1e496997",
  1216 => x"491282ca",
  1217 => x"87d8e7c0",
  1218 => x"d8d449c0",
  1219 => x"c0497487",
  1220 => x"f887e1fb",
  1221 => x"87fbf28e",
  1222 => x"711e731e",
  1223 => x"c3ff494b",
  1224 => x"fe497387",
  1225 => x"ecf287fe",
  1226 => x"1e731e87",
  1227 => x"a3c64b71",
  1228 => x"87db024a",
  1229 => x"d6028ac1",
  1230 => x"c1028a87",
  1231 => x"028a87da",
  1232 => x"8a87fcc0",
  1233 => x"87e1c002",
  1234 => x"87cb028a",
  1235 => x"c787dbc1",
  1236 => x"87c0fd49",
  1237 => x"c287dec1",
  1238 => x"02bfc4ed",
  1239 => x"4887cbc1",
  1240 => x"edc288c1",
  1241 => x"c1c158c8",
  1242 => x"c8edc287",
  1243 => x"f9c002bf",
  1244 => x"c4edc287",
  1245 => x"80c148bf",
  1246 => x"58c8edc2",
  1247 => x"c287ebc0",
  1248 => x"49bfc4ed",
  1249 => x"edc289c6",
  1250 => x"b7c059c8",
  1251 => x"87da03a9",
  1252 => x"48c4edc2",
  1253 => x"87d278c0",
  1254 => x"bfc8edc2",
  1255 => x"c287cb02",
  1256 => x"48bfc4ed",
  1257 => x"edc280c6",
  1258 => x"49c058c8",
  1259 => x"7387f6d1",
  1260 => x"fff8c049",
  1261 => x"87ddf087",
  1262 => x"5c5b5e0e",
  1263 => x"d0ff0e5d",
  1264 => x"59a6dc86",
  1265 => x"c048a6c8",
  1266 => x"c180c478",
  1267 => x"c47866c4",
  1268 => x"c478c180",
  1269 => x"c278c180",
  1270 => x"c148c8ed",
  1271 => x"ececc278",
  1272 => x"a8de48bf",
  1273 => x"f487cb05",
  1274 => x"497087db",
  1275 => x"cf59a6cc",
  1276 => x"e2e387f2",
  1277 => x"87c4e487",
  1278 => x"7087d1e3",
  1279 => x"acfbc04c",
  1280 => x"87fbc102",
  1281 => x"c10566d8",
  1282 => x"c0c187ed",
  1283 => x"82c44a66",
  1284 => x"1e727e6a",
  1285 => x"48d9e0c1",
  1286 => x"c84966c4",
  1287 => x"41204aa1",
  1288 => x"f905aa71",
  1289 => x"26511087",
  1290 => x"66c0c14a",
  1291 => x"d3c9c148",
  1292 => x"c7496a78",
  1293 => x"c1517481",
  1294 => x"c84966c0",
  1295 => x"c151c181",
  1296 => x"c94966c0",
  1297 => x"c151c081",
  1298 => x"ca4966c0",
  1299 => x"c151c081",
  1300 => x"6a1ed81e",
  1301 => x"e281c849",
  1302 => x"86c887f6",
  1303 => x"4866c4c1",
  1304 => x"c701a8c0",
  1305 => x"48a6c887",
  1306 => x"87ce78c1",
  1307 => x"4866c4c1",
  1308 => x"a6d088c1",
  1309 => x"e287c358",
  1310 => x"a6d087c2",
  1311 => x"7478c248",
  1312 => x"dbcd029c",
  1313 => x"4866c887",
  1314 => x"a866c8c1",
  1315 => x"87d0cd03",
  1316 => x"c048a6dc",
  1317 => x"c080e878",
  1318 => x"87f0e078",
  1319 => x"d0c14c70",
  1320 => x"d9c205ac",
  1321 => x"7e66c487",
  1322 => x"7087d4e3",
  1323 => x"59a6c849",
  1324 => x"7087d9e0",
  1325 => x"acecc04c",
  1326 => x"87edc105",
  1327 => x"cb4966c8",
  1328 => x"66c0c191",
  1329 => x"4aa1c481",
  1330 => x"a1c84d6a",
  1331 => x"5266c44a",
  1332 => x"79d4cac1",
  1333 => x"87f4dfff",
  1334 => x"029c4c70",
  1335 => x"fbc087d9",
  1336 => x"87d302ac",
  1337 => x"dfff5574",
  1338 => x"4c7087e2",
  1339 => x"87c7029c",
  1340 => x"05acfbc0",
  1341 => x"c087edff",
  1342 => x"c1c255e0",
  1343 => x"7d97c055",
  1344 => x"6e4966d8",
  1345 => x"87db05a9",
  1346 => x"cc4866c8",
  1347 => x"ca04a866",
  1348 => x"4866c887",
  1349 => x"a6cc80c1",
  1350 => x"cc87c858",
  1351 => x"88c14866",
  1352 => x"ff58a6d0",
  1353 => x"7087e5de",
  1354 => x"acd0c14c",
  1355 => x"d487c805",
  1356 => x"80c14866",
  1357 => x"c158a6d8",
  1358 => x"fd02acd0",
  1359 => x"e0c087e7",
  1360 => x"66d848a6",
  1361 => x"4866c478",
  1362 => x"a866e0c0",
  1363 => x"87e2c905",
  1364 => x"48a6e4c0",
  1365 => x"80c478c0",
  1366 => x"487478c0",
  1367 => x"7088fbc0",
  1368 => x"c8026e7e",
  1369 => x"486e87e5",
  1370 => x"7e7088cb",
  1371 => x"cdc1026e",
  1372 => x"c9486e87",
  1373 => x"6e7e7088",
  1374 => x"87e9c302",
  1375 => x"88c4486e",
  1376 => x"026e7e70",
  1377 => x"486e87ce",
  1378 => x"7e7088c1",
  1379 => x"d4c3026e",
  1380 => x"87f1c787",
  1381 => x"c048a6dc",
  1382 => x"dcff78f0",
  1383 => x"4c7087ee",
  1384 => x"02acecc0",
  1385 => x"c087c4c0",
  1386 => x"c05ca6e0",
  1387 => x"cd02acec",
  1388 => x"d7dcff87",
  1389 => x"c04c7087",
  1390 => x"ff05acec",
  1391 => x"ecc087f3",
  1392 => x"c4c002ac",
  1393 => x"c3dcff87",
  1394 => x"ca1ec087",
  1395 => x"4966d01e",
  1396 => x"c8c191cb",
  1397 => x"80714866",
  1398 => x"c858a6cc",
  1399 => x"80c44866",
  1400 => x"cc58a6d0",
  1401 => x"ff49bf66",
  1402 => x"c187e5dc",
  1403 => x"d41ede1e",
  1404 => x"ff49bf66",
  1405 => x"d087d9dc",
  1406 => x"c0497086",
  1407 => x"ecc08909",
  1408 => x"e8c059a6",
  1409 => x"a8c04866",
  1410 => x"87eec006",
  1411 => x"4866e8c0",
  1412 => x"c003a8dd",
  1413 => x"66c487e4",
  1414 => x"e8c049bf",
  1415 => x"e0c08166",
  1416 => x"66e8c051",
  1417 => x"c481c149",
  1418 => x"c281bf66",
  1419 => x"e8c051c1",
  1420 => x"81c24966",
  1421 => x"81bf66c4",
  1422 => x"486e51c0",
  1423 => x"78d3c9c1",
  1424 => x"81c8496e",
  1425 => x"6e5166d0",
  1426 => x"d481c949",
  1427 => x"496e5166",
  1428 => x"66dc81ca",
  1429 => x"4866d051",
  1430 => x"a6d480c1",
  1431 => x"80d84858",
  1432 => x"e6c478c1",
  1433 => x"d6dcff87",
  1434 => x"c0497087",
  1435 => x"ff59a6ec",
  1436 => x"7087ccdc",
  1437 => x"a6e0c049",
  1438 => x"4866dc59",
  1439 => x"05a8ecc0",
  1440 => x"dc87cac0",
  1441 => x"e8c048a6",
  1442 => x"c4c07866",
  1443 => x"fbd8ff87",
  1444 => x"4966c887",
  1445 => x"c0c191cb",
  1446 => x"80714866",
  1447 => x"496e7e70",
  1448 => x"4a6e81c8",
  1449 => x"e8c082ca",
  1450 => x"66dc5266",
  1451 => x"c082c14a",
  1452 => x"c18a66e8",
  1453 => x"70307248",
  1454 => x"728ac14a",
  1455 => x"69977997",
  1456 => x"ecc01e49",
  1457 => x"d9d74966",
  1458 => x"c086c487",
  1459 => x"6e58a6f0",
  1460 => x"6981c449",
  1461 => x"66e0c04d",
  1462 => x"a866c448",
  1463 => x"87c8c002",
  1464 => x"c048a6c4",
  1465 => x"87c5c078",
  1466 => x"c148a6c4",
  1467 => x"1e66c478",
  1468 => x"751ee0c0",
  1469 => x"d7d8ff49",
  1470 => x"7086c887",
  1471 => x"acb7c04c",
  1472 => x"87d4c106",
  1473 => x"e0c08574",
  1474 => x"75897449",
  1475 => x"e2e0c14b",
  1476 => x"e6fe714a",
  1477 => x"85c287d2",
  1478 => x"4866e4c0",
  1479 => x"e8c080c1",
  1480 => x"ecc058a6",
  1481 => x"81c14966",
  1482 => x"c002a970",
  1483 => x"a6c487c8",
  1484 => x"c078c048",
  1485 => x"a6c487c5",
  1486 => x"c478c148",
  1487 => x"a4c21e66",
  1488 => x"48e0c049",
  1489 => x"49708871",
  1490 => x"ff49751e",
  1491 => x"c887c1d7",
  1492 => x"a8b7c086",
  1493 => x"87c0ff01",
  1494 => x"0266e4c0",
  1495 => x"6e87d1c0",
  1496 => x"c081c949",
  1497 => x"6e5166e4",
  1498 => x"e4cbc148",
  1499 => x"87ccc078",
  1500 => x"81c9496e",
  1501 => x"486e51c2",
  1502 => x"78d8ccc1",
  1503 => x"48a6e8c0",
  1504 => x"c6c078c1",
  1505 => x"f3d5ff87",
  1506 => x"c04c7087",
  1507 => x"c00266e8",
  1508 => x"66c887f5",
  1509 => x"a866cc48",
  1510 => x"87cbc004",
  1511 => x"c14866c8",
  1512 => x"58a6cc80",
  1513 => x"cc87e0c0",
  1514 => x"88c14866",
  1515 => x"c058a6d0",
  1516 => x"c6c187d5",
  1517 => x"c8c005ac",
  1518 => x"4866d087",
  1519 => x"a6d480c1",
  1520 => x"f7d4ff58",
  1521 => x"d44c7087",
  1522 => x"80c14866",
  1523 => x"7458a6d8",
  1524 => x"cbc0029c",
  1525 => x"4866c887",
  1526 => x"a866c8c1",
  1527 => x"87f0f204",
  1528 => x"87cfd4ff",
  1529 => x"c74866c8",
  1530 => x"e5c003a8",
  1531 => x"c8edc287",
  1532 => x"c878c048",
  1533 => x"91cb4966",
  1534 => x"8166c0c1",
  1535 => x"6a4aa1c4",
  1536 => x"7952c04a",
  1537 => x"c14866c8",
  1538 => x"58a6cc80",
  1539 => x"ff04a8c7",
  1540 => x"d0ff87db",
  1541 => x"f8deff8e",
  1542 => x"616f4c87",
  1543 => x"2e2a2064",
  1544 => x"203a0020",
  1545 => x"1e731e00",
  1546 => x"029b4b71",
  1547 => x"edc287c6",
  1548 => x"78c048c4",
  1549 => x"edc21ec7",
  1550 => x"1e49bfc4",
  1551 => x"1ed4e4c1",
  1552 => x"bfececc2",
  1553 => x"87f0ed49",
  1554 => x"ecc286cc",
  1555 => x"e949bfec",
  1556 => x"9b7387ea",
  1557 => x"c187c802",
  1558 => x"c049d4e4",
  1559 => x"ff87e7e7",
  1560 => x"1e87f2dd",
  1561 => x"48c0e4c1",
  1562 => x"e5c150c0",
  1563 => x"ff49bff7",
  1564 => x"c087ead8",
  1565 => x"1e4f2648",
  1566 => x"c187e3c7",
  1567 => x"87e5fe49",
  1568 => x"87cce9fe",
  1569 => x"cd029870",
  1570 => x"c7f2fe87",
  1571 => x"02987087",
  1572 => x"4ac187c4",
  1573 => x"4ac087c2",
  1574 => x"ce059a72",
  1575 => x"c11ec087",
  1576 => x"c049c7e3",
  1577 => x"c487f7f2",
  1578 => x"c087fe86",
  1579 => x"d2e3c11e",
  1580 => x"e9f2c049",
  1581 => x"fe1ec087",
  1582 => x"497087e9",
  1583 => x"87def2c0",
  1584 => x"f887dac3",
  1585 => x"534f268e",
  1586 => x"61662044",
  1587 => x"64656c69",
  1588 => x"6f42002e",
  1589 => x"6e69746f",
  1590 => x"2e2e2e67",
  1591 => x"eac01e00",
  1592 => x"f5c087c0",
  1593 => x"87f687ee",
  1594 => x"c21e4f26",
  1595 => x"c048c4ed",
  1596 => x"ececc278",
  1597 => x"fd78c048",
  1598 => x"87e187fd",
  1599 => x"4f2648c0",
  1600 => x"00010000",
  1601 => x"20800000",
  1602 => x"74697845",
  1603 => x"42208000",
  1604 => x"006b6361",
  1605 => x"00001294",
  1606 => x"00002b58",
  1607 => x"94000000",
  1608 => x"76000012",
  1609 => x"0000002b",
  1610 => x"12940000",
  1611 => x"2b940000",
  1612 => x"00000000",
  1613 => x"00129400",
  1614 => x"002bb200",
  1615 => x"00000000",
  1616 => x"00001294",
  1617 => x"00002bd0",
  1618 => x"94000000",
  1619 => x"ee000012",
  1620 => x"0000002b",
  1621 => x"12940000",
  1622 => x"2c0c0000",
  1623 => x"00000000",
  1624 => x"00129400",
  1625 => x"00000000",
  1626 => x"00000000",
  1627 => x"00001329",
  1628 => x"00000000",
  1629 => x"7b000000",
  1630 => x"43000019",
  1631 => x"20203436",
  1632 => x"52202020",
  1633 => x"1e004d4f",
  1634 => x"c048f0fe",
  1635 => x"7909cd78",
  1636 => x"1e4f2609",
  1637 => x"bff0fe1e",
  1638 => x"2626487e",
  1639 => x"f0fe1e4f",
  1640 => x"2678c148",
  1641 => x"f0fe1e4f",
  1642 => x"2678c048",
  1643 => x"4a711e4f",
  1644 => x"265252c0",
  1645 => x"5b5e0e4f",
  1646 => x"f40e5d5c",
  1647 => x"974d7186",
  1648 => x"a5c17e6d",
  1649 => x"486c974c",
  1650 => x"6e58a6c8",
  1651 => x"a866c448",
  1652 => x"ff87c505",
  1653 => x"87e6c048",
  1654 => x"c287caff",
  1655 => x"6c9749a5",
  1656 => x"4ba3714b",
  1657 => x"974b6b97",
  1658 => x"486e7e6c",
  1659 => x"a6c880c1",
  1660 => x"cc98c758",
  1661 => x"977058a6",
  1662 => x"87e1fe7c",
  1663 => x"8ef44873",
  1664 => x"4c264d26",
  1665 => x"4f264b26",
  1666 => x"5c5b5e0e",
  1667 => x"7186f40e",
  1668 => x"4a66d84c",
  1669 => x"c29affc3",
  1670 => x"6c974ba4",
  1671 => x"49a17349",
  1672 => x"6c975172",
  1673 => x"c1486e7e",
  1674 => x"58a6c880",
  1675 => x"a6cc98c7",
  1676 => x"f4547058",
  1677 => x"87caff8e",
  1678 => x"e8fd1e1e",
  1679 => x"4abfe087",
  1680 => x"c0e0c049",
  1681 => x"87cb0299",
  1682 => x"f0c21e72",
  1683 => x"f7fe49ea",
  1684 => x"fc86c487",
  1685 => x"7e7087fd",
  1686 => x"2687c2fd",
  1687 => x"c21e4f26",
  1688 => x"fd49eaf0",
  1689 => x"e8c187c7",
  1690 => x"dafc49f8",
  1691 => x"87c7c487",
  1692 => x"ff1e4f26",
  1693 => x"e1c848d0",
  1694 => x"48d4ff78",
  1695 => x"66c478c5",
  1696 => x"c387c302",
  1697 => x"66c878e0",
  1698 => x"ff87c602",
  1699 => x"f0c348d4",
  1700 => x"48d4ff78",
  1701 => x"d0ff7871",
  1702 => x"78e1c848",
  1703 => x"2678e0c0",
  1704 => x"5b5e0e4f",
  1705 => x"4c710e5c",
  1706 => x"49eaf0c2",
  1707 => x"7087c6fc",
  1708 => x"aab7c04a",
  1709 => x"87e2c204",
  1710 => x"05aaf0c3",
  1711 => x"edc187c9",
  1712 => x"78c148e6",
  1713 => x"c387c3c2",
  1714 => x"c905aae0",
  1715 => x"eaedc187",
  1716 => x"c178c148",
  1717 => x"edc187f4",
  1718 => x"c602bfea",
  1719 => x"a2c0c287",
  1720 => x"7287c24b",
  1721 => x"059c744b",
  1722 => x"edc187d1",
  1723 => x"c11ebfe6",
  1724 => x"1ebfeaed",
  1725 => x"f9fd4972",
  1726 => x"c186c887",
  1727 => x"02bfe6ed",
  1728 => x"7387e0c0",
  1729 => x"29b7c449",
  1730 => x"c6efc191",
  1731 => x"cf4a7381",
  1732 => x"c192c29a",
  1733 => x"70307248",
  1734 => x"72baff4a",
  1735 => x"70986948",
  1736 => x"7387db79",
  1737 => x"29b7c449",
  1738 => x"c6efc191",
  1739 => x"cf4a7381",
  1740 => x"c392c29a",
  1741 => x"70307248",
  1742 => x"b069484a",
  1743 => x"edc17970",
  1744 => x"78c048ea",
  1745 => x"48e6edc1",
  1746 => x"f0c278c0",
  1747 => x"e4f949ea",
  1748 => x"c04a7087",
  1749 => x"fd03aab7",
  1750 => x"48c087de",
  1751 => x"4d2687c2",
  1752 => x"4b264c26",
  1753 => x"00004f26",
  1754 => x"00000000",
  1755 => x"711e0000",
  1756 => x"ecfc494a",
  1757 => x"1e4f2687",
  1758 => x"49724ac0",
  1759 => x"efc191c4",
  1760 => x"79c081c6",
  1761 => x"b7d082c1",
  1762 => x"87ee04aa",
  1763 => x"5e0e4f26",
  1764 => x"0e5d5c5b",
  1765 => x"ccf84d71",
  1766 => x"c44a7587",
  1767 => x"c1922ab7",
  1768 => x"7582c6ef",
  1769 => x"c29ccf4c",
  1770 => x"4b496a94",
  1771 => x"9bc32b74",
  1772 => x"307448c2",
  1773 => x"bcff4c70",
  1774 => x"98714874",
  1775 => x"dcf77a70",
  1776 => x"fe487387",
  1777 => x"000087d8",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"ff1e0000",
  1794 => x"e1c848d0",
  1795 => x"ff487178",
  1796 => x"267808d4",
  1797 => x"d0ff1e4f",
  1798 => x"78e1c848",
  1799 => x"d4ff4871",
  1800 => x"66c47808",
  1801 => x"08d4ff48",
  1802 => x"1e4f2678",
  1803 => x"66c44a71",
  1804 => x"49721e49",
  1805 => x"ff87deff",
  1806 => x"e0c048d0",
  1807 => x"4f262678",
  1808 => x"711e731e",
  1809 => x"4966c84b",
  1810 => x"c14a731e",
  1811 => x"ff49a2e0",
  1812 => x"c42687d9",
  1813 => x"264d2687",
  1814 => x"264b264c",
  1815 => x"d4ff1e4f",
  1816 => x"7affc34a",
  1817 => x"c048d0ff",
  1818 => x"7ade78e1",
  1819 => x"bff4f0c2",
  1820 => x"c848497a",
  1821 => x"717a7028",
  1822 => x"7028d048",
  1823 => x"d848717a",
  1824 => x"c27a7028",
  1825 => x"7abff8f0",
  1826 => x"28c84849",
  1827 => x"48717a70",
  1828 => x"7a7028d0",
  1829 => x"28d84871",
  1830 => x"d0ff7a70",
  1831 => x"78e0c048",
  1832 => x"731e4f26",
  1833 => x"c24a711e",
  1834 => x"4bbff4f0",
  1835 => x"e0c02b72",
  1836 => x"87ce04aa",
  1837 => x"e0c04972",
  1838 => x"f8f0c289",
  1839 => x"2b714bbf",
  1840 => x"e0c087cf",
  1841 => x"c2897249",
  1842 => x"48bff8f0",
  1843 => x"49703071",
  1844 => x"9b66c8b3",
  1845 => x"87c44873",
  1846 => x"4c264d26",
  1847 => x"4f264b26",
  1848 => x"5c5b5e0e",
  1849 => x"86ec0e5d",
  1850 => x"f0c24b71",
  1851 => x"4c7ebff4",
  1852 => x"e0c02c73",
  1853 => x"e0c004ab",
  1854 => x"48a6c487",
  1855 => x"497378c0",
  1856 => x"7189e0c0",
  1857 => x"66e4c04a",
  1858 => x"cc307248",
  1859 => x"f0c258a6",
  1860 => x"4c4dbff8",
  1861 => x"e4c02c71",
  1862 => x"c0497387",
  1863 => x"714866e4",
  1864 => x"58a6c830",
  1865 => x"7349e0c0",
  1866 => x"66e4c089",
  1867 => x"cc287148",
  1868 => x"f0c258a6",
  1869 => x"484dbff8",
  1870 => x"49703071",
  1871 => x"66e4c0b4",
  1872 => x"c084c19c",
  1873 => x"04ac66e8",
  1874 => x"4cc087c2",
  1875 => x"04abe0c0",
  1876 => x"a6cc87d3",
  1877 => x"7378c048",
  1878 => x"89e0c049",
  1879 => x"30714874",
  1880 => x"d558a6d4",
  1881 => x"74497387",
  1882 => x"d0307148",
  1883 => x"e0c058a6",
  1884 => x"74897349",
  1885 => x"d4287148",
  1886 => x"66c458a6",
  1887 => x"6ebaff4a",
  1888 => x"4966c89a",
  1889 => x"9975b9ff",
  1890 => x"66cc4872",
  1891 => x"f8f0c2b0",
  1892 => x"d0487158",
  1893 => x"f0c2b066",
  1894 => x"c0fb58fc",
  1895 => x"fc8eec87",
  1896 => x"ff1e87f6",
  1897 => x"c9c848d0",
  1898 => x"ff487178",
  1899 => x"267808d4",
  1900 => x"4a711e4f",
  1901 => x"ff87eb49",
  1902 => x"78c848d0",
  1903 => x"731e4f26",
  1904 => x"c24b711e",
  1905 => x"02bfc8f1",
  1906 => x"ebc287c3",
  1907 => x"48d0ff87",
  1908 => x"7378c9c8",
  1909 => x"b1e0c049",
  1910 => x"7148d4ff",
  1911 => x"fcf0c278",
  1912 => x"c878c048",
  1913 => x"87c50266",
  1914 => x"c249ffc3",
  1915 => x"c249c087",
  1916 => x"cc59c4f1",
  1917 => x"87c60266",
  1918 => x"4ad5d5c5",
  1919 => x"ffcf87c4",
  1920 => x"f1c24aff",
  1921 => x"f1c25ac8",
  1922 => x"78c148c8",
  1923 => x"4d2687c4",
  1924 => x"4b264c26",
  1925 => x"5e0e4f26",
  1926 => x"0e5d5c5b",
  1927 => x"f1c24a71",
  1928 => x"724cbfc4",
  1929 => x"87cb029a",
  1930 => x"c191c849",
  1931 => x"714bf4f6",
  1932 => x"c187c483",
  1933 => x"c04bf4fa",
  1934 => x"7449134d",
  1935 => x"c0f1c299",
  1936 => x"d4ffb9bf",
  1937 => x"c1787148",
  1938 => x"c8852cb7",
  1939 => x"e804adb7",
  1940 => x"fcf0c287",
  1941 => x"80c848bf",
  1942 => x"58c0f1c2",
  1943 => x"1e87effe",
  1944 => x"4b711e73",
  1945 => x"029a4a13",
  1946 => x"497287cb",
  1947 => x"1387e7fe",
  1948 => x"f5059a4a",
  1949 => x"87dafe87",
  1950 => x"fcf0c21e",
  1951 => x"f0c249bf",
  1952 => x"a1c148fc",
  1953 => x"b7c0c478",
  1954 => x"87db03a9",
  1955 => x"c248d4ff",
  1956 => x"78bfc0f1",
  1957 => x"bffcf0c2",
  1958 => x"fcf0c249",
  1959 => x"78a1c148",
  1960 => x"a9b7c0c4",
  1961 => x"ff87e504",
  1962 => x"78c848d0",
  1963 => x"48c8f1c2",
  1964 => x"4f2678c0",
  1965 => x"00000000",
  1966 => x"00000000",
  1967 => x"5f000000",
  1968 => x"0000005f",
  1969 => x"00030300",
  1970 => x"00000303",
  1971 => x"147f7f14",
  1972 => x"00147f7f",
  1973 => x"6b2e2400",
  1974 => x"00123a6b",
  1975 => x"18366a4c",
  1976 => x"0032566c",
  1977 => x"594f7e30",
  1978 => x"40683a77",
  1979 => x"07040000",
  1980 => x"00000003",
  1981 => x"3e1c0000",
  1982 => x"00004163",
  1983 => x"63410000",
  1984 => x"00001c3e",
  1985 => x"1c3e2a08",
  1986 => x"082a3e1c",
  1987 => x"3e080800",
  1988 => x"0008083e",
  1989 => x"e0800000",
  1990 => x"00000060",
  1991 => x"08080800",
  1992 => x"00080808",
  1993 => x"60000000",
  1994 => x"00000060",
  1995 => x"18306040",
  1996 => x"0103060c",
  1997 => x"597f3e00",
  1998 => x"003e7f4d",
  1999 => x"7f060400",
  2000 => x"0000007f",
  2001 => x"71634200",
  2002 => x"00464f59",
  2003 => x"49632200",
  2004 => x"00367f49",
  2005 => x"13161c18",
  2006 => x"00107f7f",
  2007 => x"45672700",
  2008 => x"00397d45",
  2009 => x"4b7e3c00",
  2010 => x"00307949",
  2011 => x"71010100",
  2012 => x"00070f79",
  2013 => x"497f3600",
  2014 => x"00367f49",
  2015 => x"494f0600",
  2016 => x"001e3f69",
  2017 => x"66000000",
  2018 => x"00000066",
  2019 => x"e6800000",
  2020 => x"00000066",
  2021 => x"14080800",
  2022 => x"00222214",
  2023 => x"14141400",
  2024 => x"00141414",
  2025 => x"14222200",
  2026 => x"00080814",
  2027 => x"51030200",
  2028 => x"00060f59",
  2029 => x"5d417f3e",
  2030 => x"001e1f55",
  2031 => x"097f7e00",
  2032 => x"007e7f09",
  2033 => x"497f7f00",
  2034 => x"00367f49",
  2035 => x"633e1c00",
  2036 => x"00414141",
  2037 => x"417f7f00",
  2038 => x"001c3e63",
  2039 => x"497f7f00",
  2040 => x"00414149",
  2041 => x"097f7f00",
  2042 => x"00010109",
  2043 => x"417f3e00",
  2044 => x"007a7b49",
  2045 => x"087f7f00",
  2046 => x"007f7f08",
  2047 => x"7f410000",
  2048 => x"0000417f",
  2049 => x"40602000",
  2050 => x"003f7f40",
  2051 => x"1c087f7f",
  2052 => x"00416336",
  2053 => x"407f7f00",
  2054 => x"00404040",
  2055 => x"0c067f7f",
  2056 => x"007f7f06",
  2057 => x"0c067f7f",
  2058 => x"007f7f18",
  2059 => x"417f3e00",
  2060 => x"003e7f41",
  2061 => x"097f7f00",
  2062 => x"00060f09",
  2063 => x"61417f3e",
  2064 => x"00407e7f",
  2065 => x"097f7f00",
  2066 => x"00667f19",
  2067 => x"4d6f2600",
  2068 => x"00327b59",
  2069 => x"7f010100",
  2070 => x"0001017f",
  2071 => x"407f3f00",
  2072 => x"003f7f40",
  2073 => x"703f0f00",
  2074 => x"000f3f70",
  2075 => x"18307f7f",
  2076 => x"007f7f30",
  2077 => x"1c366341",
  2078 => x"4163361c",
  2079 => x"7c060301",
  2080 => x"0103067c",
  2081 => x"4d597161",
  2082 => x"00414347",
  2083 => x"7f7f0000",
  2084 => x"00004141",
  2085 => x"0c060301",
  2086 => x"40603018",
  2087 => x"41410000",
  2088 => x"00007f7f",
  2089 => x"03060c08",
  2090 => x"00080c06",
  2091 => x"80808080",
  2092 => x"00808080",
  2093 => x"03000000",
  2094 => x"00000407",
  2095 => x"54742000",
  2096 => x"00787c54",
  2097 => x"447f7f00",
  2098 => x"00387c44",
  2099 => x"447c3800",
  2100 => x"00004444",
  2101 => x"447c3800",
  2102 => x"007f7f44",
  2103 => x"547c3800",
  2104 => x"00185c54",
  2105 => x"7f7e0400",
  2106 => x"00000505",
  2107 => x"a4bc1800",
  2108 => x"007cfca4",
  2109 => x"047f7f00",
  2110 => x"00787c04",
  2111 => x"3d000000",
  2112 => x"0000407d",
  2113 => x"80808000",
  2114 => x"00007dfd",
  2115 => x"107f7f00",
  2116 => x"00446c38",
  2117 => x"3f000000",
  2118 => x"0000407f",
  2119 => x"180c7c7c",
  2120 => x"00787c0c",
  2121 => x"047c7c00",
  2122 => x"00787c04",
  2123 => x"447c3800",
  2124 => x"00387c44",
  2125 => x"24fcfc00",
  2126 => x"00183c24",
  2127 => x"243c1800",
  2128 => x"00fcfc24",
  2129 => x"047c7c00",
  2130 => x"00080c04",
  2131 => x"545c4800",
  2132 => x"00207454",
  2133 => x"7f3f0400",
  2134 => x"00004444",
  2135 => x"407c3c00",
  2136 => x"007c7c40",
  2137 => x"603c1c00",
  2138 => x"001c3c60",
  2139 => x"30607c3c",
  2140 => x"003c7c60",
  2141 => x"10386c44",
  2142 => x"00446c38",
  2143 => x"e0bc1c00",
  2144 => x"001c3c60",
  2145 => x"74644400",
  2146 => x"00444c5c",
  2147 => x"3e080800",
  2148 => x"00414177",
  2149 => x"7f000000",
  2150 => x"0000007f",
  2151 => x"77414100",
  2152 => x"0008083e",
  2153 => x"03010102",
  2154 => x"00010202",
  2155 => x"7f7f7f7f",
  2156 => x"007f7f7f",
  2157 => x"1c1c0808",
  2158 => x"7f7f3e3e",
  2159 => x"3e3e7f7f",
  2160 => x"08081c1c",
  2161 => x"7c181000",
  2162 => x"0010187c",
  2163 => x"7c301000",
  2164 => x"0010307c",
  2165 => x"60603010",
  2166 => x"00061e78",
  2167 => x"183c6642",
  2168 => x"0042663c",
  2169 => x"c26a3878",
  2170 => x"00386cc6",
  2171 => x"60000060",
  2172 => x"00600000",
  2173 => x"5c5b5e0e",
  2174 => x"711e0e5d",
  2175 => x"d9f1c24c",
  2176 => x"4bc04dbf",
  2177 => x"ab741ec0",
  2178 => x"c487c702",
  2179 => x"78c048a6",
  2180 => x"a6c487c5",
  2181 => x"c478c148",
  2182 => x"49731e66",
  2183 => x"c887dfee",
  2184 => x"49e0c086",
  2185 => x"c487efef",
  2186 => x"496a4aa5",
  2187 => x"f187f0f0",
  2188 => x"85cb87c6",
  2189 => x"b7c883c1",
  2190 => x"c7ff04ab",
  2191 => x"4d262687",
  2192 => x"4b264c26",
  2193 => x"711e4f26",
  2194 => x"ddf1c24a",
  2195 => x"ddf1c25a",
  2196 => x"4978c748",
  2197 => x"2687ddfe",
  2198 => x"1e731e4f",
  2199 => x"b7c04a71",
  2200 => x"87d303aa",
  2201 => x"bff3d6c2",
  2202 => x"c187c405",
  2203 => x"c087c24b",
  2204 => x"f7d6c24b",
  2205 => x"c287c45b",
  2206 => x"c25af7d6",
  2207 => x"4abff3d6",
  2208 => x"c0c19ac1",
  2209 => x"e8ec49a2",
  2210 => x"c248fc87",
  2211 => x"78bff3d6",
  2212 => x"1e87effe",
  2213 => x"66c44a71",
  2214 => x"e649721e",
  2215 => x"262687e2",
  2216 => x"d6c21e4f",
  2217 => x"e349bff3",
  2218 => x"f1c287c4",
  2219 => x"bfe848d1",
  2220 => x"cdf1c278",
  2221 => x"78bfec48",
  2222 => x"bfd1f1c2",
  2223 => x"ffc3494a",
  2224 => x"2ab7c899",
  2225 => x"b0714872",
  2226 => x"58d9f1c2",
  2227 => x"5e0e4f26",
  2228 => x"0e5d5c5b",
  2229 => x"c8ff4b71",
  2230 => x"ccf1c287",
  2231 => x"7350c048",
  2232 => x"87eae249",
  2233 => x"c24c4970",
  2234 => x"49eecb9c",
  2235 => x"7087cccb",
  2236 => x"f1c24d49",
  2237 => x"05bf97cc",
  2238 => x"d087e2c1",
  2239 => x"f1c24966",
  2240 => x"0599bfd5",
  2241 => x"66d487d6",
  2242 => x"cdf1c249",
  2243 => x"cb0599bf",
  2244 => x"e1497387",
  2245 => x"987087f8",
  2246 => x"87c1c102",
  2247 => x"c0fe4cc1",
  2248 => x"ca497587",
  2249 => x"987087e1",
  2250 => x"c287c602",
  2251 => x"c148ccf1",
  2252 => x"ccf1c250",
  2253 => x"c005bf97",
  2254 => x"f1c287e3",
  2255 => x"d049bfd5",
  2256 => x"ff059966",
  2257 => x"f1c287d6",
  2258 => x"d449bfcd",
  2259 => x"ff059966",
  2260 => x"497387ca",
  2261 => x"7087f7e0",
  2262 => x"fffe0598",
  2263 => x"fb487487",
  2264 => x"5e0e87dc",
  2265 => x"0e5d5c5b",
  2266 => x"4dc086f4",
  2267 => x"7ebfec4c",
  2268 => x"c248a6c4",
  2269 => x"78bfd9f1",
  2270 => x"1ec01ec1",
  2271 => x"cdfd49c7",
  2272 => x"7086c887",
  2273 => x"87ce0298",
  2274 => x"ccfb49ff",
  2275 => x"49dac187",
  2276 => x"87fadfff",
  2277 => x"f1c24dc1",
  2278 => x"02bf97cc",
  2279 => x"c4d087c3",
  2280 => x"d1f1c287",
  2281 => x"d6c24bbf",
  2282 => x"c005bff3",
  2283 => x"fdc387eb",
  2284 => x"d9dfff49",
  2285 => x"49fac387",
  2286 => x"87d2dfff",
  2287 => x"ffc34973",
  2288 => x"c01e7199",
  2289 => x"87cbfb49",
  2290 => x"b7c84973",
  2291 => x"c11e7129",
  2292 => x"87fffa49",
  2293 => x"c0c686c8",
  2294 => x"d5f1c287",
  2295 => x"029b4bbf",
  2296 => x"d6c287dd",
  2297 => x"c749bfef",
  2298 => x"987087dd",
  2299 => x"c087c405",
  2300 => x"c287d24b",
  2301 => x"c2c749e0",
  2302 => x"f3d6c287",
  2303 => x"c287c658",
  2304 => x"c048efd6",
  2305 => x"c2497378",
  2306 => x"87ce0599",
  2307 => x"ff49ebc3",
  2308 => x"7087fbdd",
  2309 => x"0299c249",
  2310 => x"4cfb87c2",
  2311 => x"99c14973",
  2312 => x"c387ce05",
  2313 => x"ddff49f4",
  2314 => x"497087e4",
  2315 => x"c20299c2",
  2316 => x"734cfa87",
  2317 => x"0599c849",
  2318 => x"f5c387ce",
  2319 => x"cdddff49",
  2320 => x"c2497087",
  2321 => x"87d50299",
  2322 => x"bfddf1c2",
  2323 => x"4887ca02",
  2324 => x"f1c288c1",
  2325 => x"c2c058e1",
  2326 => x"c14cff87",
  2327 => x"c449734d",
  2328 => x"87ce0599",
  2329 => x"ff49f2c3",
  2330 => x"7087e3dc",
  2331 => x"0299c249",
  2332 => x"f1c287dc",
  2333 => x"487ebfdd",
  2334 => x"03a8b7c7",
  2335 => x"6e87cbc0",
  2336 => x"c280c148",
  2337 => x"c058e1f1",
  2338 => x"4cfe87c2",
  2339 => x"fdc34dc1",
  2340 => x"f9dbff49",
  2341 => x"c2497087",
  2342 => x"87d50299",
  2343 => x"bfddf1c2",
  2344 => x"87c9c002",
  2345 => x"48ddf1c2",
  2346 => x"c2c078c0",
  2347 => x"c14cfd87",
  2348 => x"49fac34d",
  2349 => x"87d6dbff",
  2350 => x"99c24970",
  2351 => x"87d9c002",
  2352 => x"bfddf1c2",
  2353 => x"a8b7c748",
  2354 => x"87c9c003",
  2355 => x"48ddf1c2",
  2356 => x"c2c078c7",
  2357 => x"c14cfc87",
  2358 => x"acb7c04d",
  2359 => x"87d1c003",
  2360 => x"c14a66c4",
  2361 => x"026a82d8",
  2362 => x"6a87c6c0",
  2363 => x"7349744b",
  2364 => x"c31ec00f",
  2365 => x"dac11ef0",
  2366 => x"87d2f749",
  2367 => x"987086c8",
  2368 => x"87e2c002",
  2369 => x"c248a6c8",
  2370 => x"78bfddf1",
  2371 => x"cb4966c8",
  2372 => x"4866c491",
  2373 => x"7e708071",
  2374 => x"c002bf6e",
  2375 => x"bf6e87c8",
  2376 => x"4966c84b",
  2377 => x"9d750f73",
  2378 => x"87c8c002",
  2379 => x"bfddf1c2",
  2380 => x"87c0f349",
  2381 => x"bff7d6c2",
  2382 => x"87ddc002",
  2383 => x"87c7c249",
  2384 => x"c0029870",
  2385 => x"f1c287d3",
  2386 => x"f249bfdd",
  2387 => x"49c087e6",
  2388 => x"c287c6f4",
  2389 => x"c048f7d6",
  2390 => x"f38ef478",
  2391 => x"5e0e87e0",
  2392 => x"0e5d5c5b",
  2393 => x"c24c711e",
  2394 => x"49bfd9f1",
  2395 => x"4da1cdc1",
  2396 => x"6981d1c1",
  2397 => x"029c747e",
  2398 => x"a5c487cf",
  2399 => x"c27b744b",
  2400 => x"49bfd9f1",
  2401 => x"6e87fff2",
  2402 => x"059c747b",
  2403 => x"4bc087c4",
  2404 => x"4bc187c2",
  2405 => x"c0f34973",
  2406 => x"0266d487",
  2407 => x"da4987c7",
  2408 => x"c24a7087",
  2409 => x"c24ac087",
  2410 => x"265afbd6",
  2411 => x"0087cff2",
  2412 => x"00000000",
  2413 => x"00000000",
  2414 => x"1e000000",
  2415 => x"c8ff4a71",
  2416 => x"a17249bf",
  2417 => x"1e4f2648",
  2418 => x"89bfc8ff",
  2419 => x"c0c0c0fe",
  2420 => x"01a9c0c0",
  2421 => x"4ac087c4",
  2422 => x"4ac187c2",
  2423 => x"4f264872",
  2424 => x"5c5b5e0e",
  2425 => x"4b710e5d",
  2426 => x"d04cd4ff",
  2427 => x"78c04866",
  2428 => x"d8ff49d6",
  2429 => x"ffc387d0",
  2430 => x"c3496c7c",
  2431 => x"4d7199ff",
  2432 => x"99f0c349",
  2433 => x"05a9e0c1",
  2434 => x"ffc387cb",
  2435 => x"c3486c7c",
  2436 => x"0866d098",
  2437 => x"7cffc378",
  2438 => x"c8494a6c",
  2439 => x"7cffc331",
  2440 => x"b2714a6c",
  2441 => x"31c84972",
  2442 => x"6c7cffc3",
  2443 => x"72b2714a",
  2444 => x"c331c849",
  2445 => x"4a6c7cff",
  2446 => x"d0ffb271",
  2447 => x"78e0c048",
  2448 => x"c2029b73",
  2449 => x"757b7287",
  2450 => x"264d2648",
  2451 => x"264b264c",
  2452 => x"4f261e4f",
  2453 => x"5c5b5e0e",
  2454 => x"7686f80e",
  2455 => x"49a6c81e",
  2456 => x"c487fdfd",
  2457 => x"6e4b7086",
  2458 => x"03a8c248",
  2459 => x"7387f0c2",
  2460 => x"9af0c34a",
  2461 => x"02aad0c1",
  2462 => x"e0c187c7",
  2463 => x"dec205aa",
  2464 => x"c8497387",
  2465 => x"87c30299",
  2466 => x"7387c6ff",
  2467 => x"c29cc34c",
  2468 => x"c2c105ac",
  2469 => x"4966c487",
  2470 => x"1e7131c9",
  2471 => x"d44a66c4",
  2472 => x"e1f1c292",
  2473 => x"fe817249",
  2474 => x"d887e7cc",
  2475 => x"d5d5ff49",
  2476 => x"1ec0c887",
  2477 => x"49fadfc2",
  2478 => x"87e3e8fd",
  2479 => x"c048d0ff",
  2480 => x"dfc278e0",
  2481 => x"66cc1efa",
  2482 => x"c292d44a",
  2483 => x"7249e1f1",
  2484 => x"eecafe81",
  2485 => x"c186cc87",
  2486 => x"c2c105ac",
  2487 => x"4966c487",
  2488 => x"1e7131c9",
  2489 => x"d44a66c4",
  2490 => x"e1f1c292",
  2491 => x"fe817249",
  2492 => x"c287dfcb",
  2493 => x"c81efadf",
  2494 => x"92d44a66",
  2495 => x"49e1f1c2",
  2496 => x"c8fe8172",
  2497 => x"49d787ee",
  2498 => x"87fad3ff",
  2499 => x"c21ec0c8",
  2500 => x"fd49fadf",
  2501 => x"cc87e1e6",
  2502 => x"48d0ff86",
  2503 => x"f878e0c0",
  2504 => x"87e7fc8e",
  2505 => x"5c5b5e0e",
  2506 => x"711e0e5d",
  2507 => x"4cd4ff4d",
  2508 => x"487e66d4",
  2509 => x"06a8b7c3",
  2510 => x"48c087c5",
  2511 => x"7587e2c1",
  2512 => x"f2d9fe49",
  2513 => x"c41e7587",
  2514 => x"93d44b66",
  2515 => x"83e1f1c2",
  2516 => x"c2fe4973",
  2517 => x"83c887eb",
  2518 => x"d0ff4b6b",
  2519 => x"78e1c848",
  2520 => x"49737cdd",
  2521 => x"7199ffc3",
  2522 => x"c849737c",
  2523 => x"ffc329b7",
  2524 => x"737c7199",
  2525 => x"29b7d049",
  2526 => x"7199ffc3",
  2527 => x"d849737c",
  2528 => x"7c7129b7",
  2529 => x"7c7c7cc0",
  2530 => x"7c7c7c7c",
  2531 => x"7c7c7c7c",
  2532 => x"78e0c07c",
  2533 => x"dc1e66c4",
  2534 => x"ced2ff49",
  2535 => x"7386c887",
  2536 => x"e4fa2648",
  2537 => x"dfc21e87",
  2538 => x"c149bfce",
  2539 => x"d2dfc2b9",
  2540 => x"48d4ff59",
  2541 => x"ff78ffc3",
  2542 => x"e1c048d0",
  2543 => x"48d4ff78",
  2544 => x"31c478c1",
  2545 => x"d0ff7871",
  2546 => x"78e0c048",
  2547 => x"00004f26",
  2548 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
