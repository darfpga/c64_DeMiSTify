
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"cc",x"f2",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"cc",x"f2",x"c2"),
    14 => (x"48",x"d4",x"df",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"df",x"e2"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"c4",x"4a",x"71",x"1e"),
    47 => (x"c1",x"48",x"49",x"66"),
    48 => (x"58",x"a6",x"c8",x"88"),
    49 => (x"d4",x"02",x"99",x"71"),
    50 => (x"ff",x"48",x"12",x"87"),
    51 => (x"c4",x"78",x"08",x"d4"),
    52 => (x"c1",x"48",x"49",x"66"),
    53 => (x"58",x"a6",x"c8",x"88"),
    54 => (x"ec",x"05",x"99",x"71"),
    55 => (x"1e",x"4f",x"26",x"87"),
    56 => (x"66",x"c4",x"4a",x"71"),
    57 => (x"88",x"c1",x"48",x"49"),
    58 => (x"71",x"58",x"a6",x"c8"),
    59 => (x"87",x"d6",x"02",x"99"),
    60 => (x"c3",x"48",x"d4",x"ff"),
    61 => (x"52",x"68",x"78",x"ff"),
    62 => (x"48",x"49",x"66",x"c4"),
    63 => (x"a6",x"c8",x"88",x"c1"),
    64 => (x"05",x"99",x"71",x"58"),
    65 => (x"4f",x"26",x"87",x"ea"),
    66 => (x"ff",x"1e",x"73",x"1e"),
    67 => (x"ff",x"c3",x"4b",x"d4"),
    68 => (x"c3",x"4a",x"6b",x"7b"),
    69 => (x"49",x"6b",x"7b",x"ff"),
    70 => (x"b1",x"72",x"32",x"c8"),
    71 => (x"6b",x"7b",x"ff",x"c3"),
    72 => (x"71",x"31",x"c8",x"4a"),
    73 => (x"7b",x"ff",x"c3",x"b2"),
    74 => (x"32",x"c8",x"49",x"6b"),
    75 => (x"48",x"71",x"b1",x"72"),
    76 => (x"4d",x"26",x"87",x"c4"),
    77 => (x"4b",x"26",x"4c",x"26"),
    78 => (x"5e",x"0e",x"4f",x"26"),
    79 => (x"0e",x"5d",x"5c",x"5b"),
    80 => (x"d4",x"ff",x"4a",x"71"),
    81 => (x"c3",x"49",x"72",x"4c"),
    82 => (x"7c",x"71",x"99",x"ff"),
    83 => (x"bf",x"d4",x"df",x"c2"),
    84 => (x"d0",x"87",x"c8",x"05"),
    85 => (x"30",x"c9",x"48",x"66"),
    86 => (x"d0",x"58",x"a6",x"d4"),
    87 => (x"29",x"d8",x"49",x"66"),
    88 => (x"71",x"99",x"ff",x"c3"),
    89 => (x"49",x"66",x"d0",x"7c"),
    90 => (x"ff",x"c3",x"29",x"d0"),
    91 => (x"d0",x"7c",x"71",x"99"),
    92 => (x"29",x"c8",x"49",x"66"),
    93 => (x"71",x"99",x"ff",x"c3"),
    94 => (x"49",x"66",x"d0",x"7c"),
    95 => (x"71",x"99",x"ff",x"c3"),
    96 => (x"d0",x"49",x"72",x"7c"),
    97 => (x"99",x"ff",x"c3",x"29"),
    98 => (x"4b",x"6c",x"7c",x"71"),
    99 => (x"4d",x"ff",x"f0",x"c9"),
   100 => (x"05",x"ab",x"ff",x"c3"),
   101 => (x"ff",x"c3",x"87",x"d0"),
   102 => (x"c1",x"4b",x"6c",x"7c"),
   103 => (x"87",x"c6",x"02",x"8d"),
   104 => (x"02",x"ab",x"ff",x"c3"),
   105 => (x"48",x"73",x"87",x"f0"),
   106 => (x"1e",x"87",x"c7",x"fe"),
   107 => (x"d4",x"ff",x"49",x"c0"),
   108 => (x"78",x"ff",x"c3",x"48"),
   109 => (x"c8",x"c3",x"81",x"c1"),
   110 => (x"f1",x"04",x"a9",x"b7"),
   111 => (x"1e",x"4f",x"26",x"87"),
   112 => (x"87",x"e7",x"1e",x"73"),
   113 => (x"4b",x"df",x"f8",x"c4"),
   114 => (x"ff",x"c0",x"1e",x"c0"),
   115 => (x"49",x"f7",x"c1",x"f0"),
   116 => (x"c4",x"87",x"e7",x"fd"),
   117 => (x"05",x"a8",x"c1",x"86"),
   118 => (x"ff",x"87",x"ea",x"c0"),
   119 => (x"ff",x"c3",x"48",x"d4"),
   120 => (x"c0",x"c0",x"c1",x"78"),
   121 => (x"1e",x"c0",x"c0",x"c0"),
   122 => (x"c1",x"f0",x"e1",x"c0"),
   123 => (x"c9",x"fd",x"49",x"e9"),
   124 => (x"70",x"86",x"c4",x"87"),
   125 => (x"87",x"ca",x"05",x"98"),
   126 => (x"c3",x"48",x"d4",x"ff"),
   127 => (x"48",x"c1",x"78",x"ff"),
   128 => (x"e6",x"fe",x"87",x"cb"),
   129 => (x"05",x"8b",x"c1",x"87"),
   130 => (x"c0",x"87",x"fd",x"fe"),
   131 => (x"87",x"e6",x"fc",x"48"),
   132 => (x"ff",x"1e",x"73",x"1e"),
   133 => (x"ff",x"c3",x"48",x"d4"),
   134 => (x"c0",x"4b",x"d3",x"78"),
   135 => (x"f0",x"ff",x"c0",x"1e"),
   136 => (x"fc",x"49",x"c1",x"c1"),
   137 => (x"86",x"c4",x"87",x"d4"),
   138 => (x"ca",x"05",x"98",x"70"),
   139 => (x"48",x"d4",x"ff",x"87"),
   140 => (x"c1",x"78",x"ff",x"c3"),
   141 => (x"fd",x"87",x"cb",x"48"),
   142 => (x"8b",x"c1",x"87",x"f1"),
   143 => (x"87",x"db",x"ff",x"05"),
   144 => (x"f1",x"fb",x"48",x"c0"),
   145 => (x"5b",x"5e",x"0e",x"87"),
   146 => (x"d4",x"ff",x"0e",x"5c"),
   147 => (x"87",x"db",x"fd",x"4c"),
   148 => (x"c0",x"1e",x"ea",x"c6"),
   149 => (x"c8",x"c1",x"f0",x"e1"),
   150 => (x"87",x"de",x"fb",x"49"),
   151 => (x"a8",x"c1",x"86",x"c4"),
   152 => (x"fe",x"87",x"c8",x"02"),
   153 => (x"48",x"c0",x"87",x"ea"),
   154 => (x"fa",x"87",x"e2",x"c1"),
   155 => (x"49",x"70",x"87",x"da"),
   156 => (x"99",x"ff",x"ff",x"cf"),
   157 => (x"02",x"a9",x"ea",x"c6"),
   158 => (x"d3",x"fe",x"87",x"c8"),
   159 => (x"c1",x"48",x"c0",x"87"),
   160 => (x"ff",x"c3",x"87",x"cb"),
   161 => (x"4b",x"f1",x"c0",x"7c"),
   162 => (x"70",x"87",x"f4",x"fc"),
   163 => (x"eb",x"c0",x"02",x"98"),
   164 => (x"c0",x"1e",x"c0",x"87"),
   165 => (x"fa",x"c1",x"f0",x"ff"),
   166 => (x"87",x"de",x"fa",x"49"),
   167 => (x"98",x"70",x"86",x"c4"),
   168 => (x"c3",x"87",x"d9",x"05"),
   169 => (x"49",x"6c",x"7c",x"ff"),
   170 => (x"7c",x"7c",x"ff",x"c3"),
   171 => (x"c0",x"c1",x"7c",x"7c"),
   172 => (x"87",x"c4",x"02",x"99"),
   173 => (x"87",x"d5",x"48",x"c1"),
   174 => (x"87",x"d1",x"48",x"c0"),
   175 => (x"c4",x"05",x"ab",x"c2"),
   176 => (x"c8",x"48",x"c0",x"87"),
   177 => (x"05",x"8b",x"c1",x"87"),
   178 => (x"c0",x"87",x"fd",x"fe"),
   179 => (x"87",x"e4",x"f9",x"48"),
   180 => (x"c2",x"1e",x"73",x"1e"),
   181 => (x"c1",x"48",x"d4",x"df"),
   182 => (x"ff",x"4b",x"c7",x"78"),
   183 => (x"78",x"c2",x"48",x"d0"),
   184 => (x"ff",x"87",x"c8",x"fb"),
   185 => (x"78",x"c3",x"48",x"d0"),
   186 => (x"e5",x"c0",x"1e",x"c0"),
   187 => (x"49",x"c0",x"c1",x"d0"),
   188 => (x"c4",x"87",x"c7",x"f9"),
   189 => (x"05",x"a8",x"c1",x"86"),
   190 => (x"c2",x"4b",x"87",x"c1"),
   191 => (x"87",x"c5",x"05",x"ab"),
   192 => (x"f9",x"c0",x"48",x"c0"),
   193 => (x"05",x"8b",x"c1",x"87"),
   194 => (x"fc",x"87",x"d0",x"ff"),
   195 => (x"df",x"c2",x"87",x"f7"),
   196 => (x"98",x"70",x"58",x"d8"),
   197 => (x"c1",x"87",x"cd",x"05"),
   198 => (x"f0",x"ff",x"c0",x"1e"),
   199 => (x"f8",x"49",x"d0",x"c1"),
   200 => (x"86",x"c4",x"87",x"d8"),
   201 => (x"c3",x"48",x"d4",x"ff"),
   202 => (x"de",x"c4",x"78",x"ff"),
   203 => (x"dc",x"df",x"c2",x"87"),
   204 => (x"48",x"d0",x"ff",x"58"),
   205 => (x"d4",x"ff",x"78",x"c2"),
   206 => (x"78",x"ff",x"c3",x"48"),
   207 => (x"f5",x"f7",x"48",x"c1"),
   208 => (x"5b",x"5e",x"0e",x"87"),
   209 => (x"71",x"0e",x"5d",x"5c"),
   210 => (x"4d",x"ff",x"c3",x"4a"),
   211 => (x"75",x"4c",x"d4",x"ff"),
   212 => (x"48",x"d0",x"ff",x"7c"),
   213 => (x"75",x"78",x"c3",x"c4"),
   214 => (x"c0",x"1e",x"72",x"7c"),
   215 => (x"d8",x"c1",x"f0",x"ff"),
   216 => (x"87",x"d6",x"f7",x"49"),
   217 => (x"98",x"70",x"86",x"c4"),
   218 => (x"c1",x"87",x"c5",x"02"),
   219 => (x"87",x"f0",x"c0",x"48"),
   220 => (x"fe",x"c3",x"7c",x"75"),
   221 => (x"1e",x"c0",x"c8",x"7c"),
   222 => (x"f4",x"49",x"66",x"d4"),
   223 => (x"86",x"c4",x"87",x"fa"),
   224 => (x"7c",x"75",x"7c",x"75"),
   225 => (x"da",x"d8",x"7c",x"75"),
   226 => (x"7c",x"75",x"4b",x"e0"),
   227 => (x"05",x"99",x"49",x"6c"),
   228 => (x"8b",x"c1",x"87",x"c5"),
   229 => (x"75",x"87",x"f3",x"05"),
   230 => (x"48",x"d0",x"ff",x"7c"),
   231 => (x"48",x"c0",x"78",x"c2"),
   232 => (x"0e",x"87",x"cf",x"f6"),
   233 => (x"5d",x"5c",x"5b",x"5e"),
   234 => (x"c0",x"4b",x"71",x"0e"),
   235 => (x"cd",x"ee",x"c5",x"4c"),
   236 => (x"d4",x"ff",x"4a",x"df"),
   237 => (x"78",x"ff",x"c3",x"48"),
   238 => (x"fe",x"c3",x"49",x"68"),
   239 => (x"fd",x"c0",x"05",x"a9"),
   240 => (x"73",x"4d",x"70",x"87"),
   241 => (x"87",x"cc",x"02",x"9b"),
   242 => (x"73",x"1e",x"66",x"d0"),
   243 => (x"87",x"cf",x"f4",x"49"),
   244 => (x"87",x"d6",x"86",x"c4"),
   245 => (x"c4",x"48",x"d0",x"ff"),
   246 => (x"ff",x"c3",x"78",x"d1"),
   247 => (x"48",x"66",x"d0",x"7d"),
   248 => (x"a6",x"d4",x"88",x"c1"),
   249 => (x"05",x"98",x"70",x"58"),
   250 => (x"d4",x"ff",x"87",x"f0"),
   251 => (x"78",x"ff",x"c3",x"48"),
   252 => (x"05",x"9b",x"73",x"78"),
   253 => (x"d0",x"ff",x"87",x"c5"),
   254 => (x"c1",x"78",x"d0",x"48"),
   255 => (x"8a",x"c1",x"4c",x"4a"),
   256 => (x"87",x"ee",x"fe",x"05"),
   257 => (x"e9",x"f4",x"48",x"74"),
   258 => (x"1e",x"73",x"1e",x"87"),
   259 => (x"4b",x"c0",x"4a",x"71"),
   260 => (x"c3",x"48",x"d4",x"ff"),
   261 => (x"d0",x"ff",x"78",x"ff"),
   262 => (x"78",x"c3",x"c4",x"48"),
   263 => (x"c3",x"48",x"d4",x"ff"),
   264 => (x"1e",x"72",x"78",x"ff"),
   265 => (x"c1",x"f0",x"ff",x"c0"),
   266 => (x"cd",x"f4",x"49",x"d1"),
   267 => (x"70",x"86",x"c4",x"87"),
   268 => (x"87",x"d2",x"05",x"98"),
   269 => (x"cc",x"1e",x"c0",x"c8"),
   270 => (x"e6",x"fd",x"49",x"66"),
   271 => (x"70",x"86",x"c4",x"87"),
   272 => (x"48",x"d0",x"ff",x"4b"),
   273 => (x"48",x"73",x"78",x"c2"),
   274 => (x"0e",x"87",x"eb",x"f3"),
   275 => (x"5d",x"5c",x"5b",x"5e"),
   276 => (x"c0",x"1e",x"c0",x"0e"),
   277 => (x"c9",x"c1",x"f0",x"ff"),
   278 => (x"87",x"de",x"f3",x"49"),
   279 => (x"df",x"c2",x"1e",x"d2"),
   280 => (x"fe",x"fc",x"49",x"dc"),
   281 => (x"c0",x"86",x"c8",x"87"),
   282 => (x"d2",x"84",x"c1",x"4c"),
   283 => (x"f8",x"04",x"ac",x"b7"),
   284 => (x"dc",x"df",x"c2",x"87"),
   285 => (x"c3",x"49",x"bf",x"97"),
   286 => (x"c0",x"c1",x"99",x"c0"),
   287 => (x"e7",x"c0",x"05",x"a9"),
   288 => (x"e3",x"df",x"c2",x"87"),
   289 => (x"d0",x"49",x"bf",x"97"),
   290 => (x"e4",x"df",x"c2",x"31"),
   291 => (x"c8",x"4a",x"bf",x"97"),
   292 => (x"c2",x"b1",x"72",x"32"),
   293 => (x"bf",x"97",x"e5",x"df"),
   294 => (x"4c",x"71",x"b1",x"4a"),
   295 => (x"ff",x"ff",x"ff",x"cf"),
   296 => (x"ca",x"84",x"c1",x"9c"),
   297 => (x"87",x"e7",x"c1",x"34"),
   298 => (x"97",x"e5",x"df",x"c2"),
   299 => (x"31",x"c1",x"49",x"bf"),
   300 => (x"df",x"c2",x"99",x"c6"),
   301 => (x"4a",x"bf",x"97",x"e6"),
   302 => (x"72",x"2a",x"b7",x"c7"),
   303 => (x"e1",x"df",x"c2",x"b1"),
   304 => (x"4d",x"4a",x"bf",x"97"),
   305 => (x"df",x"c2",x"9d",x"cf"),
   306 => (x"4a",x"bf",x"97",x"e2"),
   307 => (x"32",x"ca",x"9a",x"c3"),
   308 => (x"97",x"e3",x"df",x"c2"),
   309 => (x"33",x"c2",x"4b",x"bf"),
   310 => (x"df",x"c2",x"b2",x"73"),
   311 => (x"4b",x"bf",x"97",x"e4"),
   312 => (x"c6",x"9b",x"c0",x"c3"),
   313 => (x"b2",x"73",x"2b",x"b7"),
   314 => (x"48",x"c1",x"81",x"c2"),
   315 => (x"49",x"70",x"30",x"71"),
   316 => (x"30",x"75",x"48",x"c1"),
   317 => (x"4c",x"72",x"4d",x"70"),
   318 => (x"94",x"71",x"84",x"c1"),
   319 => (x"ad",x"b7",x"c0",x"c8"),
   320 => (x"c1",x"87",x"cc",x"06"),
   321 => (x"c8",x"2d",x"b7",x"34"),
   322 => (x"01",x"ad",x"b7",x"c0"),
   323 => (x"74",x"87",x"f4",x"ff"),
   324 => (x"87",x"de",x"f0",x"48"),
   325 => (x"5c",x"5b",x"5e",x"0e"),
   326 => (x"86",x"f8",x"0e",x"5d"),
   327 => (x"48",x"c2",x"e8",x"c2"),
   328 => (x"df",x"c2",x"78",x"c0"),
   329 => (x"49",x"c0",x"1e",x"fa"),
   330 => (x"c4",x"87",x"de",x"fb"),
   331 => (x"05",x"98",x"70",x"86"),
   332 => (x"48",x"c0",x"87",x"c5"),
   333 => (x"c0",x"87",x"ce",x"c9"),
   334 => (x"c0",x"7e",x"c1",x"4d"),
   335 => (x"49",x"bf",x"f6",x"f2"),
   336 => (x"4a",x"f0",x"e0",x"c2"),
   337 => (x"ec",x"4b",x"c8",x"71"),
   338 => (x"98",x"70",x"87",x"e0"),
   339 => (x"c0",x"87",x"c2",x"05"),
   340 => (x"f2",x"f2",x"c0",x"7e"),
   341 => (x"e1",x"c2",x"49",x"bf"),
   342 => (x"c8",x"71",x"4a",x"cc"),
   343 => (x"87",x"ca",x"ec",x"4b"),
   344 => (x"c2",x"05",x"98",x"70"),
   345 => (x"6e",x"7e",x"c0",x"87"),
   346 => (x"87",x"fd",x"c0",x"02"),
   347 => (x"bf",x"c0",x"e7",x"c2"),
   348 => (x"f8",x"e7",x"c2",x"4d"),
   349 => (x"48",x"7e",x"bf",x"9f"),
   350 => (x"a8",x"ea",x"d6",x"c5"),
   351 => (x"c2",x"87",x"c7",x"05"),
   352 => (x"4d",x"bf",x"c0",x"e7"),
   353 => (x"48",x"6e",x"87",x"ce"),
   354 => (x"a8",x"d5",x"e9",x"ca"),
   355 => (x"c0",x"87",x"c5",x"02"),
   356 => (x"87",x"f1",x"c7",x"48"),
   357 => (x"1e",x"fa",x"df",x"c2"),
   358 => (x"ec",x"f9",x"49",x"75"),
   359 => (x"70",x"86",x"c4",x"87"),
   360 => (x"87",x"c5",x"05",x"98"),
   361 => (x"dc",x"c7",x"48",x"c0"),
   362 => (x"f2",x"f2",x"c0",x"87"),
   363 => (x"e1",x"c2",x"49",x"bf"),
   364 => (x"c8",x"71",x"4a",x"cc"),
   365 => (x"87",x"f2",x"ea",x"4b"),
   366 => (x"c8",x"05",x"98",x"70"),
   367 => (x"c2",x"e8",x"c2",x"87"),
   368 => (x"da",x"78",x"c1",x"48"),
   369 => (x"f6",x"f2",x"c0",x"87"),
   370 => (x"e0",x"c2",x"49",x"bf"),
   371 => (x"c8",x"71",x"4a",x"f0"),
   372 => (x"87",x"d6",x"ea",x"4b"),
   373 => (x"c0",x"02",x"98",x"70"),
   374 => (x"48",x"c0",x"87",x"c5"),
   375 => (x"c2",x"87",x"e6",x"c6"),
   376 => (x"bf",x"97",x"f8",x"e7"),
   377 => (x"a9",x"d5",x"c1",x"49"),
   378 => (x"87",x"cd",x"c0",x"05"),
   379 => (x"97",x"f9",x"e7",x"c2"),
   380 => (x"ea",x"c2",x"49",x"bf"),
   381 => (x"c5",x"c0",x"02",x"a9"),
   382 => (x"c6",x"48",x"c0",x"87"),
   383 => (x"df",x"c2",x"87",x"c7"),
   384 => (x"7e",x"bf",x"97",x"fa"),
   385 => (x"a8",x"e9",x"c3",x"48"),
   386 => (x"87",x"ce",x"c0",x"02"),
   387 => (x"eb",x"c3",x"48",x"6e"),
   388 => (x"c5",x"c0",x"02",x"a8"),
   389 => (x"c5",x"48",x"c0",x"87"),
   390 => (x"e0",x"c2",x"87",x"eb"),
   391 => (x"49",x"bf",x"97",x"c5"),
   392 => (x"cc",x"c0",x"05",x"99"),
   393 => (x"c6",x"e0",x"c2",x"87"),
   394 => (x"c2",x"49",x"bf",x"97"),
   395 => (x"c5",x"c0",x"02",x"a9"),
   396 => (x"c5",x"48",x"c0",x"87"),
   397 => (x"e0",x"c2",x"87",x"cf"),
   398 => (x"48",x"bf",x"97",x"c7"),
   399 => (x"58",x"fe",x"e7",x"c2"),
   400 => (x"c1",x"48",x"4c",x"70"),
   401 => (x"c2",x"e8",x"c2",x"88"),
   402 => (x"c8",x"e0",x"c2",x"58"),
   403 => (x"75",x"49",x"bf",x"97"),
   404 => (x"c9",x"e0",x"c2",x"81"),
   405 => (x"c8",x"4a",x"bf",x"97"),
   406 => (x"7e",x"a1",x"72",x"32"),
   407 => (x"48",x"cf",x"ec",x"c2"),
   408 => (x"e0",x"c2",x"78",x"6e"),
   409 => (x"48",x"bf",x"97",x"ca"),
   410 => (x"c2",x"58",x"a6",x"c8"),
   411 => (x"02",x"bf",x"c2",x"e8"),
   412 => (x"c0",x"87",x"d4",x"c2"),
   413 => (x"49",x"bf",x"f2",x"f2"),
   414 => (x"4a",x"cc",x"e1",x"c2"),
   415 => (x"e7",x"4b",x"c8",x"71"),
   416 => (x"98",x"70",x"87",x"e8"),
   417 => (x"87",x"c5",x"c0",x"02"),
   418 => (x"f8",x"c3",x"48",x"c0"),
   419 => (x"fa",x"e7",x"c2",x"87"),
   420 => (x"ec",x"c2",x"4c",x"bf"),
   421 => (x"e0",x"c2",x"5c",x"e3"),
   422 => (x"49",x"bf",x"97",x"df"),
   423 => (x"e0",x"c2",x"31",x"c8"),
   424 => (x"4a",x"bf",x"97",x"de"),
   425 => (x"e0",x"c2",x"49",x"a1"),
   426 => (x"4a",x"bf",x"97",x"e0"),
   427 => (x"a1",x"72",x"32",x"d0"),
   428 => (x"e1",x"e0",x"c2",x"49"),
   429 => (x"d8",x"4a",x"bf",x"97"),
   430 => (x"49",x"a1",x"72",x"32"),
   431 => (x"c2",x"91",x"66",x"c4"),
   432 => (x"81",x"bf",x"cf",x"ec"),
   433 => (x"59",x"d7",x"ec",x"c2"),
   434 => (x"97",x"e7",x"e0",x"c2"),
   435 => (x"32",x"c8",x"4a",x"bf"),
   436 => (x"97",x"e6",x"e0",x"c2"),
   437 => (x"4a",x"a2",x"4b",x"bf"),
   438 => (x"97",x"e8",x"e0",x"c2"),
   439 => (x"33",x"d0",x"4b",x"bf"),
   440 => (x"c2",x"4a",x"a2",x"73"),
   441 => (x"bf",x"97",x"e9",x"e0"),
   442 => (x"d8",x"9b",x"cf",x"4b"),
   443 => (x"4a",x"a2",x"73",x"33"),
   444 => (x"5a",x"db",x"ec",x"c2"),
   445 => (x"bf",x"d7",x"ec",x"c2"),
   446 => (x"74",x"8a",x"c2",x"4a"),
   447 => (x"db",x"ec",x"c2",x"92"),
   448 => (x"78",x"a1",x"72",x"48"),
   449 => (x"c2",x"87",x"ca",x"c1"),
   450 => (x"bf",x"97",x"cc",x"e0"),
   451 => (x"c2",x"31",x"c8",x"49"),
   452 => (x"bf",x"97",x"cb",x"e0"),
   453 => (x"c2",x"49",x"a1",x"4a"),
   454 => (x"c2",x"59",x"ca",x"e8"),
   455 => (x"49",x"bf",x"c6",x"e8"),
   456 => (x"ff",x"c7",x"31",x"c5"),
   457 => (x"c2",x"29",x"c9",x"81"),
   458 => (x"c2",x"59",x"e3",x"ec"),
   459 => (x"bf",x"97",x"d1",x"e0"),
   460 => (x"c2",x"32",x"c8",x"4a"),
   461 => (x"bf",x"97",x"d0",x"e0"),
   462 => (x"c4",x"4a",x"a2",x"4b"),
   463 => (x"82",x"6e",x"92",x"66"),
   464 => (x"5a",x"df",x"ec",x"c2"),
   465 => (x"48",x"d7",x"ec",x"c2"),
   466 => (x"ec",x"c2",x"78",x"c0"),
   467 => (x"a1",x"72",x"48",x"d3"),
   468 => (x"e3",x"ec",x"c2",x"78"),
   469 => (x"d7",x"ec",x"c2",x"48"),
   470 => (x"ec",x"c2",x"78",x"bf"),
   471 => (x"ec",x"c2",x"48",x"e7"),
   472 => (x"c2",x"78",x"bf",x"db"),
   473 => (x"02",x"bf",x"c2",x"e8"),
   474 => (x"74",x"87",x"c9",x"c0"),
   475 => (x"70",x"30",x"c4",x"48"),
   476 => (x"87",x"c9",x"c0",x"7e"),
   477 => (x"bf",x"df",x"ec",x"c2"),
   478 => (x"70",x"30",x"c4",x"48"),
   479 => (x"c6",x"e8",x"c2",x"7e"),
   480 => (x"c1",x"78",x"6e",x"48"),
   481 => (x"26",x"8e",x"f8",x"48"),
   482 => (x"26",x"4c",x"26",x"4d"),
   483 => (x"0e",x"4f",x"26",x"4b"),
   484 => (x"5d",x"5c",x"5b",x"5e"),
   485 => (x"c2",x"4a",x"71",x"0e"),
   486 => (x"02",x"bf",x"c2",x"e8"),
   487 => (x"4b",x"72",x"87",x"cb"),
   488 => (x"4c",x"72",x"2b",x"c7"),
   489 => (x"c9",x"9c",x"ff",x"c1"),
   490 => (x"c8",x"4b",x"72",x"87"),
   491 => (x"c3",x"4c",x"72",x"2b"),
   492 => (x"ec",x"c2",x"9c",x"ff"),
   493 => (x"c0",x"83",x"bf",x"cf"),
   494 => (x"ab",x"bf",x"ee",x"f2"),
   495 => (x"c0",x"87",x"d9",x"02"),
   496 => (x"c2",x"5b",x"f2",x"f2"),
   497 => (x"73",x"1e",x"fa",x"df"),
   498 => (x"87",x"fd",x"f0",x"49"),
   499 => (x"98",x"70",x"86",x"c4"),
   500 => (x"c0",x"87",x"c5",x"05"),
   501 => (x"87",x"e6",x"c0",x"48"),
   502 => (x"bf",x"c2",x"e8",x"c2"),
   503 => (x"74",x"87",x"d2",x"02"),
   504 => (x"c2",x"91",x"c4",x"49"),
   505 => (x"69",x"81",x"fa",x"df"),
   506 => (x"ff",x"ff",x"cf",x"4d"),
   507 => (x"cb",x"9d",x"ff",x"ff"),
   508 => (x"c2",x"49",x"74",x"87"),
   509 => (x"fa",x"df",x"c2",x"91"),
   510 => (x"4d",x"69",x"9f",x"81"),
   511 => (x"c6",x"fe",x"48",x"75"),
   512 => (x"5b",x"5e",x"0e",x"87"),
   513 => (x"f8",x"0e",x"5d",x"5c"),
   514 => (x"9c",x"4c",x"71",x"86"),
   515 => (x"c0",x"87",x"c5",x"05"),
   516 => (x"87",x"c1",x"c3",x"48"),
   517 => (x"6e",x"7e",x"a4",x"c8"),
   518 => (x"d8",x"78",x"c0",x"48"),
   519 => (x"87",x"c7",x"02",x"66"),
   520 => (x"bf",x"97",x"66",x"d8"),
   521 => (x"c0",x"87",x"c5",x"05"),
   522 => (x"87",x"e9",x"c2",x"48"),
   523 => (x"49",x"c1",x"1e",x"c0"),
   524 => (x"c4",x"87",x"e0",x"ca"),
   525 => (x"9d",x"4d",x"70",x"86"),
   526 => (x"87",x"c2",x"c1",x"02"),
   527 => (x"4a",x"ca",x"e8",x"c2"),
   528 => (x"e0",x"49",x"66",x"d8"),
   529 => (x"98",x"70",x"87",x"c9"),
   530 => (x"87",x"f2",x"c0",x"02"),
   531 => (x"66",x"d8",x"4a",x"75"),
   532 => (x"e0",x"4b",x"cb",x"49"),
   533 => (x"98",x"70",x"87",x"ee"),
   534 => (x"87",x"e2",x"c0",x"02"),
   535 => (x"9d",x"75",x"1e",x"c0"),
   536 => (x"c8",x"87",x"c7",x"02"),
   537 => (x"78",x"c0",x"48",x"a6"),
   538 => (x"a6",x"c8",x"87",x"c5"),
   539 => (x"c8",x"78",x"c1",x"48"),
   540 => (x"de",x"c9",x"49",x"66"),
   541 => (x"70",x"86",x"c4",x"87"),
   542 => (x"fe",x"05",x"9d",x"4d"),
   543 => (x"9d",x"75",x"87",x"fe"),
   544 => (x"87",x"cf",x"c1",x"02"),
   545 => (x"6e",x"49",x"a5",x"dc"),
   546 => (x"da",x"78",x"69",x"48"),
   547 => (x"a6",x"c4",x"49",x"a5"),
   548 => (x"78",x"a4",x"c4",x"48"),
   549 => (x"c4",x"48",x"69",x"9f"),
   550 => (x"c2",x"78",x"08",x"66"),
   551 => (x"02",x"bf",x"c2",x"e8"),
   552 => (x"a5",x"d4",x"87",x"d2"),
   553 => (x"49",x"69",x"9f",x"49"),
   554 => (x"99",x"ff",x"ff",x"c0"),
   555 => (x"30",x"d0",x"48",x"71"),
   556 => (x"87",x"c2",x"7e",x"70"),
   557 => (x"49",x"6e",x"7e",x"c0"),
   558 => (x"bf",x"66",x"c4",x"48"),
   559 => (x"08",x"66",x"c4",x"80"),
   560 => (x"cc",x"7c",x"c0",x"78"),
   561 => (x"66",x"c4",x"49",x"a4"),
   562 => (x"a4",x"d0",x"79",x"bf"),
   563 => (x"c1",x"79",x"c0",x"49"),
   564 => (x"c0",x"87",x"c2",x"48"),
   565 => (x"fa",x"8e",x"f8",x"48"),
   566 => (x"5e",x"0e",x"87",x"ed"),
   567 => (x"0e",x"5d",x"5c",x"5b"),
   568 => (x"02",x"9c",x"4c",x"71"),
   569 => (x"c8",x"87",x"ca",x"c1"),
   570 => (x"02",x"69",x"49",x"a4"),
   571 => (x"d0",x"87",x"c2",x"c1"),
   572 => (x"49",x"6c",x"4a",x"66"),
   573 => (x"5a",x"a6",x"d4",x"82"),
   574 => (x"b9",x"4d",x"66",x"d0"),
   575 => (x"bf",x"fe",x"e7",x"c2"),
   576 => (x"72",x"ba",x"ff",x"4a"),
   577 => (x"02",x"99",x"71",x"99"),
   578 => (x"c4",x"87",x"e4",x"c0"),
   579 => (x"49",x"6b",x"4b",x"a4"),
   580 => (x"70",x"87",x"fc",x"f9"),
   581 => (x"fa",x"e7",x"c2",x"7b"),
   582 => (x"81",x"6c",x"49",x"bf"),
   583 => (x"b9",x"75",x"7c",x"71"),
   584 => (x"bf",x"fe",x"e7",x"c2"),
   585 => (x"72",x"ba",x"ff",x"4a"),
   586 => (x"05",x"99",x"71",x"99"),
   587 => (x"75",x"87",x"dc",x"ff"),
   588 => (x"87",x"d3",x"f9",x"7c"),
   589 => (x"71",x"1e",x"73",x"1e"),
   590 => (x"c7",x"02",x"9b",x"4b"),
   591 => (x"49",x"a3",x"c8",x"87"),
   592 => (x"87",x"c5",x"05",x"69"),
   593 => (x"f7",x"c0",x"48",x"c0"),
   594 => (x"d3",x"ec",x"c2",x"87"),
   595 => (x"a3",x"c4",x"4a",x"bf"),
   596 => (x"c2",x"49",x"69",x"49"),
   597 => (x"fa",x"e7",x"c2",x"89"),
   598 => (x"a2",x"71",x"91",x"bf"),
   599 => (x"fe",x"e7",x"c2",x"4a"),
   600 => (x"99",x"6b",x"49",x"bf"),
   601 => (x"c0",x"4a",x"a2",x"71"),
   602 => (x"c8",x"5a",x"f2",x"f2"),
   603 => (x"49",x"72",x"1e",x"66"),
   604 => (x"c4",x"87",x"d6",x"ea"),
   605 => (x"05",x"98",x"70",x"86"),
   606 => (x"48",x"c0",x"87",x"c4"),
   607 => (x"48",x"c1",x"87",x"c2"),
   608 => (x"1e",x"87",x"c8",x"f8"),
   609 => (x"4b",x"71",x"1e",x"73"),
   610 => (x"87",x"c7",x"02",x"9b"),
   611 => (x"69",x"49",x"a3",x"c8"),
   612 => (x"c0",x"87",x"c5",x"05"),
   613 => (x"87",x"f7",x"c0",x"48"),
   614 => (x"bf",x"d3",x"ec",x"c2"),
   615 => (x"49",x"a3",x"c4",x"4a"),
   616 => (x"89",x"c2",x"49",x"69"),
   617 => (x"bf",x"fa",x"e7",x"c2"),
   618 => (x"4a",x"a2",x"71",x"91"),
   619 => (x"bf",x"fe",x"e7",x"c2"),
   620 => (x"71",x"99",x"6b",x"49"),
   621 => (x"f2",x"c0",x"4a",x"a2"),
   622 => (x"66",x"c8",x"5a",x"f2"),
   623 => (x"e5",x"49",x"72",x"1e"),
   624 => (x"86",x"c4",x"87",x"ff"),
   625 => (x"c4",x"05",x"98",x"70"),
   626 => (x"c2",x"48",x"c0",x"87"),
   627 => (x"f6",x"48",x"c1",x"87"),
   628 => (x"5e",x"0e",x"87",x"f9"),
   629 => (x"1e",x"0e",x"5c",x"5b"),
   630 => (x"66",x"d0",x"4b",x"71"),
   631 => (x"73",x"2c",x"c9",x"4c"),
   632 => (x"d4",x"c1",x"02",x"9b"),
   633 => (x"49",x"a3",x"c8",x"87"),
   634 => (x"cc",x"c1",x"02",x"69"),
   635 => (x"fe",x"e7",x"c2",x"87"),
   636 => (x"b9",x"ff",x"49",x"bf"),
   637 => (x"7e",x"99",x"4a",x"6b"),
   638 => (x"d1",x"03",x"ac",x"71"),
   639 => (x"d0",x"7b",x"c0",x"87"),
   640 => (x"79",x"c0",x"49",x"a3"),
   641 => (x"c4",x"4a",x"a3",x"cc"),
   642 => (x"79",x"6a",x"49",x"a3"),
   643 => (x"8c",x"72",x"87",x"c2"),
   644 => (x"c0",x"02",x"9c",x"74"),
   645 => (x"1e",x"49",x"87",x"e3"),
   646 => (x"fd",x"fa",x"49",x"73"),
   647 => (x"d0",x"86",x"c4",x"87"),
   648 => (x"ff",x"c7",x"49",x"66"),
   649 => (x"87",x"cb",x"02",x"99"),
   650 => (x"1e",x"fa",x"df",x"c2"),
   651 => (x"c3",x"fc",x"49",x"73"),
   652 => (x"d0",x"86",x"c4",x"87"),
   653 => (x"66",x"d0",x"49",x"a3"),
   654 => (x"cc",x"f5",x"26",x"79"),
   655 => (x"1e",x"73",x"1e",x"87"),
   656 => (x"02",x"9b",x"4b",x"71"),
   657 => (x"c2",x"87",x"e4",x"c0"),
   658 => (x"73",x"5b",x"e7",x"ec"),
   659 => (x"c2",x"8a",x"c2",x"4a"),
   660 => (x"49",x"bf",x"fa",x"e7"),
   661 => (x"d3",x"ec",x"c2",x"92"),
   662 => (x"80",x"72",x"48",x"bf"),
   663 => (x"58",x"eb",x"ec",x"c2"),
   664 => (x"30",x"c4",x"48",x"71"),
   665 => (x"58",x"ca",x"e8",x"c2"),
   666 => (x"c2",x"87",x"ed",x"c0"),
   667 => (x"c2",x"48",x"e3",x"ec"),
   668 => (x"78",x"bf",x"d7",x"ec"),
   669 => (x"48",x"e7",x"ec",x"c2"),
   670 => (x"bf",x"db",x"ec",x"c2"),
   671 => (x"c2",x"e8",x"c2",x"78"),
   672 => (x"87",x"c9",x"02",x"bf"),
   673 => (x"bf",x"fa",x"e7",x"c2"),
   674 => (x"c7",x"31",x"c4",x"49"),
   675 => (x"df",x"ec",x"c2",x"87"),
   676 => (x"31",x"c4",x"49",x"bf"),
   677 => (x"59",x"ca",x"e8",x"c2"),
   678 => (x"0e",x"87",x"f0",x"f3"),
   679 => (x"0e",x"5c",x"5b",x"5e"),
   680 => (x"4b",x"c0",x"4a",x"71"),
   681 => (x"c0",x"02",x"9a",x"72"),
   682 => (x"a2",x"da",x"87",x"e1"),
   683 => (x"4b",x"69",x"9f",x"49"),
   684 => (x"bf",x"c2",x"e8",x"c2"),
   685 => (x"d4",x"87",x"cf",x"02"),
   686 => (x"69",x"9f",x"49",x"a2"),
   687 => (x"ff",x"c0",x"4c",x"49"),
   688 => (x"34",x"d0",x"9c",x"ff"),
   689 => (x"4c",x"c0",x"87",x"c2"),
   690 => (x"73",x"b3",x"49",x"74"),
   691 => (x"87",x"ed",x"fd",x"49"),
   692 => (x"0e",x"87",x"f6",x"f2"),
   693 => (x"5d",x"5c",x"5b",x"5e"),
   694 => (x"71",x"86",x"f4",x"0e"),
   695 => (x"72",x"7e",x"c0",x"4a"),
   696 => (x"87",x"d8",x"02",x"9a"),
   697 => (x"48",x"f6",x"df",x"c2"),
   698 => (x"df",x"c2",x"78",x"c0"),
   699 => (x"ec",x"c2",x"48",x"ee"),
   700 => (x"c2",x"78",x"bf",x"e7"),
   701 => (x"c2",x"48",x"f2",x"df"),
   702 => (x"78",x"bf",x"e3",x"ec"),
   703 => (x"48",x"d7",x"e8",x"c2"),
   704 => (x"e8",x"c2",x"50",x"c0"),
   705 => (x"c2",x"49",x"bf",x"c6"),
   706 => (x"4a",x"bf",x"f6",x"df"),
   707 => (x"c4",x"03",x"aa",x"71"),
   708 => (x"49",x"72",x"87",x"c9"),
   709 => (x"c0",x"05",x"99",x"cf"),
   710 => (x"f2",x"c0",x"87",x"e9"),
   711 => (x"df",x"c2",x"48",x"ee"),
   712 => (x"c2",x"78",x"bf",x"ee"),
   713 => (x"c2",x"1e",x"fa",x"df"),
   714 => (x"49",x"bf",x"ee",x"df"),
   715 => (x"48",x"ee",x"df",x"c2"),
   716 => (x"71",x"78",x"a1",x"c1"),
   717 => (x"c4",x"87",x"d2",x"e3"),
   718 => (x"ea",x"f2",x"c0",x"86"),
   719 => (x"fa",x"df",x"c2",x"48"),
   720 => (x"c0",x"87",x"cc",x"78"),
   721 => (x"48",x"bf",x"ea",x"f2"),
   722 => (x"c0",x"80",x"e0",x"c0"),
   723 => (x"c2",x"58",x"ee",x"f2"),
   724 => (x"48",x"bf",x"f6",x"df"),
   725 => (x"df",x"c2",x"80",x"c1"),
   726 => (x"aa",x"27",x"58",x"fa"),
   727 => (x"bf",x"00",x"00",x"0c"),
   728 => (x"9d",x"4d",x"bf",x"97"),
   729 => (x"87",x"e3",x"c2",x"02"),
   730 => (x"02",x"ad",x"e5",x"c3"),
   731 => (x"c0",x"87",x"dc",x"c2"),
   732 => (x"4b",x"bf",x"ea",x"f2"),
   733 => (x"11",x"49",x"a3",x"cb"),
   734 => (x"05",x"ac",x"cf",x"4c"),
   735 => (x"75",x"87",x"d2",x"c1"),
   736 => (x"c1",x"99",x"df",x"49"),
   737 => (x"c2",x"91",x"cd",x"89"),
   738 => (x"c1",x"81",x"ca",x"e8"),
   739 => (x"51",x"12",x"4a",x"a3"),
   740 => (x"12",x"4a",x"a3",x"c3"),
   741 => (x"4a",x"a3",x"c5",x"51"),
   742 => (x"a3",x"c7",x"51",x"12"),
   743 => (x"c9",x"51",x"12",x"4a"),
   744 => (x"51",x"12",x"4a",x"a3"),
   745 => (x"12",x"4a",x"a3",x"ce"),
   746 => (x"4a",x"a3",x"d0",x"51"),
   747 => (x"a3",x"d2",x"51",x"12"),
   748 => (x"d4",x"51",x"12",x"4a"),
   749 => (x"51",x"12",x"4a",x"a3"),
   750 => (x"12",x"4a",x"a3",x"d6"),
   751 => (x"4a",x"a3",x"d8",x"51"),
   752 => (x"a3",x"dc",x"51",x"12"),
   753 => (x"de",x"51",x"12",x"4a"),
   754 => (x"51",x"12",x"4a",x"a3"),
   755 => (x"fa",x"c0",x"7e",x"c1"),
   756 => (x"c8",x"49",x"74",x"87"),
   757 => (x"eb",x"c0",x"05",x"99"),
   758 => (x"d0",x"49",x"74",x"87"),
   759 => (x"87",x"d1",x"05",x"99"),
   760 => (x"c0",x"02",x"66",x"dc"),
   761 => (x"49",x"73",x"87",x"cb"),
   762 => (x"70",x"0f",x"66",x"dc"),
   763 => (x"d3",x"c0",x"02",x"98"),
   764 => (x"c0",x"05",x"6e",x"87"),
   765 => (x"e8",x"c2",x"87",x"c6"),
   766 => (x"50",x"c0",x"48",x"ca"),
   767 => (x"bf",x"ea",x"f2",x"c0"),
   768 => (x"87",x"e1",x"c2",x"48"),
   769 => (x"48",x"d7",x"e8",x"c2"),
   770 => (x"c2",x"7e",x"50",x"c0"),
   771 => (x"49",x"bf",x"c6",x"e8"),
   772 => (x"bf",x"f6",x"df",x"c2"),
   773 => (x"04",x"aa",x"71",x"4a"),
   774 => (x"c2",x"87",x"f7",x"fb"),
   775 => (x"05",x"bf",x"e7",x"ec"),
   776 => (x"c2",x"87",x"c8",x"c0"),
   777 => (x"02",x"bf",x"c2",x"e8"),
   778 => (x"c2",x"87",x"f8",x"c1"),
   779 => (x"49",x"bf",x"f2",x"df"),
   780 => (x"70",x"87",x"dc",x"ed"),
   781 => (x"f6",x"df",x"c2",x"49"),
   782 => (x"48",x"a6",x"c4",x"59"),
   783 => (x"bf",x"f2",x"df",x"c2"),
   784 => (x"c2",x"e8",x"c2",x"78"),
   785 => (x"d8",x"c0",x"02",x"bf"),
   786 => (x"49",x"66",x"c4",x"87"),
   787 => (x"ff",x"ff",x"ff",x"cf"),
   788 => (x"02",x"a9",x"99",x"f8"),
   789 => (x"c0",x"87",x"c5",x"c0"),
   790 => (x"87",x"e1",x"c0",x"4c"),
   791 => (x"dc",x"c0",x"4c",x"c1"),
   792 => (x"49",x"66",x"c4",x"87"),
   793 => (x"99",x"f8",x"ff",x"cf"),
   794 => (x"c8",x"c0",x"02",x"a9"),
   795 => (x"48",x"a6",x"c8",x"87"),
   796 => (x"c5",x"c0",x"78",x"c0"),
   797 => (x"48",x"a6",x"c8",x"87"),
   798 => (x"66",x"c8",x"78",x"c1"),
   799 => (x"05",x"9c",x"74",x"4c"),
   800 => (x"c4",x"87",x"e0",x"c0"),
   801 => (x"89",x"c2",x"49",x"66"),
   802 => (x"bf",x"fa",x"e7",x"c2"),
   803 => (x"ec",x"c2",x"91",x"4a"),
   804 => (x"c2",x"4a",x"bf",x"d3"),
   805 => (x"72",x"48",x"ee",x"df"),
   806 => (x"df",x"c2",x"78",x"a1"),
   807 => (x"78",x"c0",x"48",x"f6"),
   808 => (x"c0",x"87",x"df",x"f9"),
   809 => (x"eb",x"8e",x"f4",x"48"),
   810 => (x"00",x"00",x"87",x"dd"),
   811 => (x"ff",x"ff",x"00",x"00"),
   812 => (x"0c",x"ba",x"ff",x"ff"),
   813 => (x"0c",x"c3",x"00",x"00"),
   814 => (x"41",x"46",x"00",x"00"),
   815 => (x"20",x"32",x"33",x"54"),
   816 => (x"46",x"00",x"20",x"20"),
   817 => (x"36",x"31",x"54",x"41"),
   818 => (x"00",x"20",x"20",x"20"),
   819 => (x"48",x"d4",x"ff",x"1e"),
   820 => (x"68",x"78",x"ff",x"c3"),
   821 => (x"1e",x"4f",x"26",x"48"),
   822 => (x"c3",x"48",x"d4",x"ff"),
   823 => (x"d0",x"ff",x"78",x"ff"),
   824 => (x"78",x"e1",x"c0",x"48"),
   825 => (x"d4",x"48",x"d4",x"ff"),
   826 => (x"eb",x"ec",x"c2",x"78"),
   827 => (x"bf",x"d4",x"ff",x"48"),
   828 => (x"1e",x"4f",x"26",x"50"),
   829 => (x"c0",x"48",x"d0",x"ff"),
   830 => (x"4f",x"26",x"78",x"e0"),
   831 => (x"87",x"cc",x"ff",x"1e"),
   832 => (x"02",x"99",x"49",x"70"),
   833 => (x"fb",x"c0",x"87",x"c6"),
   834 => (x"87",x"f1",x"05",x"a9"),
   835 => (x"4f",x"26",x"48",x"71"),
   836 => (x"5c",x"5b",x"5e",x"0e"),
   837 => (x"c0",x"4b",x"71",x"0e"),
   838 => (x"87",x"f0",x"fe",x"4c"),
   839 => (x"02",x"99",x"49",x"70"),
   840 => (x"c0",x"87",x"f9",x"c0"),
   841 => (x"c0",x"02",x"a9",x"ec"),
   842 => (x"fb",x"c0",x"87",x"f2"),
   843 => (x"eb",x"c0",x"02",x"a9"),
   844 => (x"b7",x"66",x"cc",x"87"),
   845 => (x"87",x"c7",x"03",x"ac"),
   846 => (x"c2",x"02",x"66",x"d0"),
   847 => (x"71",x"53",x"71",x"87"),
   848 => (x"87",x"c2",x"02",x"99"),
   849 => (x"c3",x"fe",x"84",x"c1"),
   850 => (x"99",x"49",x"70",x"87"),
   851 => (x"c0",x"87",x"cd",x"02"),
   852 => (x"c7",x"02",x"a9",x"ec"),
   853 => (x"a9",x"fb",x"c0",x"87"),
   854 => (x"87",x"d5",x"ff",x"05"),
   855 => (x"c3",x"02",x"66",x"d0"),
   856 => (x"7b",x"97",x"c0",x"87"),
   857 => (x"05",x"a9",x"ec",x"c0"),
   858 => (x"4a",x"74",x"87",x"c4"),
   859 => (x"4a",x"74",x"87",x"c5"),
   860 => (x"72",x"8a",x"0a",x"c0"),
   861 => (x"26",x"87",x"c2",x"48"),
   862 => (x"26",x"4c",x"26",x"4d"),
   863 => (x"1e",x"4f",x"26",x"4b"),
   864 => (x"70",x"87",x"c9",x"fd"),
   865 => (x"f0",x"c0",x"4a",x"49"),
   866 => (x"87",x"c9",x"04",x"aa"),
   867 => (x"01",x"aa",x"f9",x"c0"),
   868 => (x"f0",x"c0",x"87",x"c3"),
   869 => (x"aa",x"c1",x"c1",x"8a"),
   870 => (x"c1",x"87",x"c9",x"04"),
   871 => (x"c3",x"01",x"aa",x"da"),
   872 => (x"8a",x"f7",x"c0",x"87"),
   873 => (x"04",x"aa",x"e1",x"c1"),
   874 => (x"fa",x"c1",x"87",x"c9"),
   875 => (x"87",x"c3",x"01",x"aa"),
   876 => (x"72",x"8a",x"fd",x"c0"),
   877 => (x"0e",x"4f",x"26",x"48"),
   878 => (x"0e",x"5c",x"5b",x"5e"),
   879 => (x"d4",x"ff",x"4a",x"71"),
   880 => (x"c0",x"49",x"72",x"4c"),
   881 => (x"4b",x"70",x"87",x"e9"),
   882 => (x"87",x"c2",x"02",x"9b"),
   883 => (x"d0",x"ff",x"8b",x"c1"),
   884 => (x"c1",x"78",x"c5",x"48"),
   885 => (x"49",x"73",x"7c",x"d5"),
   886 => (x"e4",x"c1",x"31",x"c6"),
   887 => (x"4a",x"bf",x"97",x"c0"),
   888 => (x"70",x"b0",x"71",x"48"),
   889 => (x"48",x"d0",x"ff",x"7c"),
   890 => (x"48",x"73",x"78",x"c4"),
   891 => (x"0e",x"87",x"ca",x"fe"),
   892 => (x"5d",x"5c",x"5b",x"5e"),
   893 => (x"71",x"86",x"f8",x"0e"),
   894 => (x"fb",x"7e",x"c0",x"4c"),
   895 => (x"4b",x"c0",x"87",x"d9"),
   896 => (x"97",x"dc",x"fa",x"c0"),
   897 => (x"a9",x"c0",x"49",x"bf"),
   898 => (x"fb",x"87",x"cf",x"04"),
   899 => (x"83",x"c1",x"87",x"ee"),
   900 => (x"97",x"dc",x"fa",x"c0"),
   901 => (x"06",x"ab",x"49",x"bf"),
   902 => (x"fa",x"c0",x"87",x"f1"),
   903 => (x"02",x"bf",x"97",x"dc"),
   904 => (x"e7",x"fa",x"87",x"cf"),
   905 => (x"99",x"49",x"70",x"87"),
   906 => (x"c0",x"87",x"c6",x"02"),
   907 => (x"f1",x"05",x"a9",x"ec"),
   908 => (x"fa",x"4b",x"c0",x"87"),
   909 => (x"4d",x"70",x"87",x"d6"),
   910 => (x"c8",x"87",x"d1",x"fa"),
   911 => (x"cb",x"fa",x"58",x"a6"),
   912 => (x"c1",x"4a",x"70",x"87"),
   913 => (x"49",x"a4",x"c8",x"83"),
   914 => (x"ad",x"49",x"69",x"97"),
   915 => (x"c0",x"87",x"c7",x"02"),
   916 => (x"c0",x"05",x"ad",x"ff"),
   917 => (x"a4",x"c9",x"87",x"e7"),
   918 => (x"49",x"69",x"97",x"49"),
   919 => (x"02",x"a9",x"66",x"c4"),
   920 => (x"c0",x"48",x"87",x"c7"),
   921 => (x"d4",x"05",x"a8",x"ff"),
   922 => (x"49",x"a4",x"ca",x"87"),
   923 => (x"aa",x"49",x"69",x"97"),
   924 => (x"c0",x"87",x"c6",x"02"),
   925 => (x"c4",x"05",x"aa",x"ff"),
   926 => (x"d0",x"7e",x"c1",x"87"),
   927 => (x"ad",x"ec",x"c0",x"87"),
   928 => (x"c0",x"87",x"c6",x"02"),
   929 => (x"c4",x"05",x"ad",x"fb"),
   930 => (x"c1",x"4b",x"c0",x"87"),
   931 => (x"fe",x"02",x"6e",x"7e"),
   932 => (x"de",x"f9",x"87",x"e1"),
   933 => (x"f8",x"48",x"73",x"87"),
   934 => (x"87",x"db",x"fb",x"8e"),
   935 => (x"5b",x"5e",x"0e",x"00"),
   936 => (x"f8",x"0e",x"5d",x"5c"),
   937 => (x"ff",x"4d",x"71",x"86"),
   938 => (x"1e",x"75",x"4b",x"d4"),
   939 => (x"49",x"f0",x"ec",x"c2"),
   940 => (x"c4",x"87",x"ce",x"e5"),
   941 => (x"02",x"98",x"70",x"86"),
   942 => (x"c4",x"87",x"d2",x"c4"),
   943 => (x"e4",x"c1",x"48",x"a6"),
   944 => (x"75",x"78",x"bf",x"c2"),
   945 => (x"87",x"ef",x"fb",x"49"),
   946 => (x"c5",x"48",x"d0",x"ff"),
   947 => (x"7b",x"d6",x"c1",x"78"),
   948 => (x"a2",x"75",x"4a",x"c0"),
   949 => (x"c1",x"7b",x"11",x"49"),
   950 => (x"aa",x"b7",x"cb",x"82"),
   951 => (x"cc",x"87",x"f3",x"04"),
   952 => (x"7b",x"ff",x"c3",x"4a"),
   953 => (x"e0",x"c0",x"82",x"c1"),
   954 => (x"f4",x"04",x"aa",x"b7"),
   955 => (x"48",x"d0",x"ff",x"87"),
   956 => (x"ff",x"c3",x"78",x"c4"),
   957 => (x"c1",x"78",x"c5",x"7b"),
   958 => (x"7b",x"c1",x"7b",x"d3"),
   959 => (x"48",x"66",x"78",x"c4"),
   960 => (x"06",x"a8",x"b7",x"c0"),
   961 => (x"c2",x"87",x"f6",x"c2"),
   962 => (x"4c",x"bf",x"f8",x"ec"),
   963 => (x"74",x"48",x"66",x"c4"),
   964 => (x"58",x"a6",x"c8",x"88"),
   965 => (x"c1",x"02",x"9c",x"74"),
   966 => (x"df",x"c2",x"87",x"ff"),
   967 => (x"c0",x"c8",x"7e",x"fa"),
   968 => (x"b7",x"c0",x"8c",x"4d"),
   969 => (x"87",x"c6",x"03",x"ac"),
   970 => (x"4d",x"a4",x"c0",x"c8"),
   971 => (x"c0",x"c8",x"4c",x"c0"),
   972 => (x"87",x"dc",x"05",x"ad"),
   973 => (x"97",x"eb",x"ec",x"c2"),
   974 => (x"99",x"d0",x"49",x"bf"),
   975 => (x"c0",x"87",x"d1",x"02"),
   976 => (x"f0",x"ec",x"c2",x"1e"),
   977 => (x"87",x"ec",x"e7",x"49"),
   978 => (x"49",x"70",x"86",x"c4"),
   979 => (x"87",x"ee",x"c0",x"4a"),
   980 => (x"1e",x"fa",x"df",x"c2"),
   981 => (x"49",x"f0",x"ec",x"c2"),
   982 => (x"c4",x"87",x"d9",x"e7"),
   983 => (x"4a",x"49",x"70",x"86"),
   984 => (x"c8",x"48",x"d0",x"ff"),
   985 => (x"d4",x"c1",x"78",x"c5"),
   986 => (x"bf",x"97",x"6e",x"7b"),
   987 => (x"c1",x"48",x"6e",x"7b"),
   988 => (x"c1",x"7e",x"70",x"80"),
   989 => (x"f0",x"ff",x"05",x"8d"),
   990 => (x"48",x"d0",x"ff",x"87"),
   991 => (x"9a",x"72",x"78",x"c4"),
   992 => (x"c0",x"87",x"c5",x"05"),
   993 => (x"87",x"c7",x"c1",x"48"),
   994 => (x"ec",x"c2",x"1e",x"c1"),
   995 => (x"c9",x"e5",x"49",x"f0"),
   996 => (x"74",x"86",x"c4",x"87"),
   997 => (x"c1",x"fe",x"05",x"9c"),
   998 => (x"48",x"66",x"c4",x"87"),
   999 => (x"06",x"a8",x"b7",x"c0"),
  1000 => (x"ec",x"c2",x"87",x"d1"),
  1001 => (x"78",x"c0",x"48",x"f0"),
  1002 => (x"78",x"c0",x"80",x"d0"),
  1003 => (x"ec",x"c2",x"80",x"f4"),
  1004 => (x"c4",x"78",x"bf",x"fc"),
  1005 => (x"b7",x"c0",x"48",x"66"),
  1006 => (x"ca",x"fd",x"01",x"a8"),
  1007 => (x"48",x"d0",x"ff",x"87"),
  1008 => (x"d3",x"c1",x"78",x"c5"),
  1009 => (x"c4",x"7b",x"c0",x"7b"),
  1010 => (x"c2",x"48",x"c1",x"78"),
  1011 => (x"f8",x"48",x"c0",x"87"),
  1012 => (x"26",x"4d",x"26",x"8e"),
  1013 => (x"26",x"4b",x"26",x"4c"),
  1014 => (x"5b",x"5e",x"0e",x"4f"),
  1015 => (x"1e",x"0e",x"5d",x"5c"),
  1016 => (x"4c",x"c0",x"4b",x"71"),
  1017 => (x"c0",x"04",x"ab",x"4d"),
  1018 => (x"f7",x"c0",x"87",x"e8"),
  1019 => (x"9d",x"75",x"1e",x"ef"),
  1020 => (x"c0",x"87",x"c4",x"02"),
  1021 => (x"c1",x"87",x"c2",x"4a"),
  1022 => (x"eb",x"49",x"72",x"4a"),
  1023 => (x"86",x"c4",x"87",x"d5"),
  1024 => (x"84",x"c1",x"7e",x"70"),
  1025 => (x"87",x"c2",x"05",x"6e"),
  1026 => (x"85",x"c1",x"4c",x"73"),
  1027 => (x"ff",x"06",x"ac",x"73"),
  1028 => (x"48",x"6e",x"87",x"d8"),
  1029 => (x"87",x"f9",x"fe",x"26"),
  1030 => (x"5c",x"5b",x"5e",x"0e"),
  1031 => (x"cc",x"4b",x"71",x"0e"),
  1032 => (x"87",x"d8",x"02",x"66"),
  1033 => (x"8c",x"f0",x"c0",x"4c"),
  1034 => (x"74",x"87",x"d8",x"02"),
  1035 => (x"02",x"8a",x"c1",x"4a"),
  1036 => (x"02",x"8a",x"87",x"d1"),
  1037 => (x"02",x"8a",x"87",x"cd"),
  1038 => (x"87",x"d9",x"87",x"c9"),
  1039 => (x"dc",x"f9",x"49",x"73"),
  1040 => (x"74",x"87",x"d2",x"87"),
  1041 => (x"c1",x"49",x"c0",x"1e"),
  1042 => (x"74",x"87",x"d9",x"db"),
  1043 => (x"c1",x"49",x"73",x"1e"),
  1044 => (x"c8",x"87",x"d1",x"db"),
  1045 => (x"87",x"fb",x"fd",x"86"),
  1046 => (x"5c",x"5b",x"5e",x"0e"),
  1047 => (x"71",x"1e",x"0e",x"5d"),
  1048 => (x"91",x"de",x"49",x"4c"),
  1049 => (x"4d",x"d8",x"ed",x"c2"),
  1050 => (x"6d",x"97",x"85",x"71"),
  1051 => (x"87",x"dc",x"c1",x"02"),
  1052 => (x"bf",x"c4",x"ed",x"c2"),
  1053 => (x"72",x"82",x"74",x"4a"),
  1054 => (x"87",x"dd",x"fd",x"49"),
  1055 => (x"02",x"6e",x"7e",x"70"),
  1056 => (x"c2",x"87",x"f2",x"c0"),
  1057 => (x"6e",x"4b",x"cc",x"ed"),
  1058 => (x"ff",x"49",x"cb",x"4a"),
  1059 => (x"74",x"87",x"d9",x"c0"),
  1060 => (x"c1",x"93",x"cb",x"4b"),
  1061 => (x"c4",x"83",x"d4",x"e4"),
  1062 => (x"d0",x"c3",x"c1",x"83"),
  1063 => (x"c1",x"49",x"74",x"7b"),
  1064 => (x"75",x"87",x"d1",x"c5"),
  1065 => (x"c1",x"e4",x"c1",x"7b"),
  1066 => (x"1e",x"49",x"bf",x"97"),
  1067 => (x"49",x"cc",x"ed",x"c2"),
  1068 => (x"c4",x"87",x"e5",x"fd"),
  1069 => (x"c1",x"49",x"74",x"86"),
  1070 => (x"c0",x"87",x"f9",x"c4"),
  1071 => (x"d8",x"c6",x"c1",x"49"),
  1072 => (x"ec",x"ec",x"c2",x"87"),
  1073 => (x"c1",x"78",x"c0",x"48"),
  1074 => (x"87",x"d9",x"dd",x"49"),
  1075 => (x"87",x"c1",x"fc",x"26"),
  1076 => (x"64",x"61",x"6f",x"4c"),
  1077 => (x"2e",x"67",x"6e",x"69"),
  1078 => (x"0e",x"00",x"2e",x"2e"),
  1079 => (x"0e",x"5c",x"5b",x"5e"),
  1080 => (x"c2",x"4a",x"4b",x"71"),
  1081 => (x"82",x"bf",x"c4",x"ed"),
  1082 => (x"ec",x"fb",x"49",x"72"),
  1083 => (x"9c",x"4c",x"70",x"87"),
  1084 => (x"49",x"87",x"c4",x"02"),
  1085 => (x"c2",x"87",x"e4",x"e6"),
  1086 => (x"c0",x"48",x"c4",x"ed"),
  1087 => (x"dc",x"49",x"c1",x"78"),
  1088 => (x"ce",x"fb",x"87",x"e3"),
  1089 => (x"5b",x"5e",x"0e",x"87"),
  1090 => (x"f4",x"0e",x"5d",x"5c"),
  1091 => (x"fa",x"df",x"c2",x"86"),
  1092 => (x"c4",x"4c",x"c0",x"4d"),
  1093 => (x"78",x"c0",x"48",x"a6"),
  1094 => (x"bf",x"c4",x"ed",x"c2"),
  1095 => (x"06",x"a9",x"c0",x"49"),
  1096 => (x"c2",x"87",x"c1",x"c1"),
  1097 => (x"98",x"48",x"fa",x"df"),
  1098 => (x"87",x"f8",x"c0",x"02"),
  1099 => (x"1e",x"ef",x"f7",x"c0"),
  1100 => (x"c7",x"02",x"66",x"c8"),
  1101 => (x"48",x"a6",x"c4",x"87"),
  1102 => (x"87",x"c5",x"78",x"c0"),
  1103 => (x"c1",x"48",x"a6",x"c4"),
  1104 => (x"49",x"66",x"c4",x"78"),
  1105 => (x"c4",x"87",x"cc",x"e6"),
  1106 => (x"c1",x"4d",x"70",x"86"),
  1107 => (x"48",x"66",x"c4",x"84"),
  1108 => (x"a6",x"c8",x"80",x"c1"),
  1109 => (x"c4",x"ed",x"c2",x"58"),
  1110 => (x"03",x"ac",x"49",x"bf"),
  1111 => (x"9d",x"75",x"87",x"c6"),
  1112 => (x"87",x"c8",x"ff",x"05"),
  1113 => (x"9d",x"75",x"4c",x"c0"),
  1114 => (x"87",x"e0",x"c3",x"02"),
  1115 => (x"1e",x"ef",x"f7",x"c0"),
  1116 => (x"c7",x"02",x"66",x"c8"),
  1117 => (x"48",x"a6",x"cc",x"87"),
  1118 => (x"87",x"c5",x"78",x"c0"),
  1119 => (x"c1",x"48",x"a6",x"cc"),
  1120 => (x"49",x"66",x"cc",x"78"),
  1121 => (x"c4",x"87",x"cc",x"e5"),
  1122 => (x"6e",x"7e",x"70",x"86"),
  1123 => (x"87",x"e9",x"c2",x"02"),
  1124 => (x"81",x"cb",x"49",x"6e"),
  1125 => (x"d0",x"49",x"69",x"97"),
  1126 => (x"d6",x"c1",x"02",x"99"),
  1127 => (x"db",x"c3",x"c1",x"87"),
  1128 => (x"cb",x"49",x"74",x"4a"),
  1129 => (x"d4",x"e4",x"c1",x"91"),
  1130 => (x"c8",x"79",x"72",x"81"),
  1131 => (x"51",x"ff",x"c3",x"81"),
  1132 => (x"91",x"de",x"49",x"74"),
  1133 => (x"4d",x"d8",x"ed",x"c2"),
  1134 => (x"c1",x"c2",x"85",x"71"),
  1135 => (x"a5",x"c1",x"7d",x"97"),
  1136 => (x"51",x"e0",x"c0",x"49"),
  1137 => (x"97",x"ca",x"e8",x"c2"),
  1138 => (x"87",x"d2",x"02",x"bf"),
  1139 => (x"a5",x"c2",x"84",x"c1"),
  1140 => (x"ca",x"e8",x"c2",x"4b"),
  1141 => (x"fe",x"49",x"db",x"4a"),
  1142 => (x"c1",x"87",x"cd",x"fb"),
  1143 => (x"a5",x"cd",x"87",x"db"),
  1144 => (x"c1",x"51",x"c0",x"49"),
  1145 => (x"4b",x"a5",x"c2",x"84"),
  1146 => (x"49",x"cb",x"4a",x"6e"),
  1147 => (x"87",x"f8",x"fa",x"fe"),
  1148 => (x"c1",x"87",x"c6",x"c1"),
  1149 => (x"74",x"4a",x"d8",x"c1"),
  1150 => (x"c1",x"91",x"cb",x"49"),
  1151 => (x"72",x"81",x"d4",x"e4"),
  1152 => (x"ca",x"e8",x"c2",x"79"),
  1153 => (x"d8",x"02",x"bf",x"97"),
  1154 => (x"de",x"49",x"74",x"87"),
  1155 => (x"c2",x"84",x"c1",x"91"),
  1156 => (x"71",x"4b",x"d8",x"ed"),
  1157 => (x"ca",x"e8",x"c2",x"83"),
  1158 => (x"fe",x"49",x"dd",x"4a"),
  1159 => (x"d8",x"87",x"c9",x"fa"),
  1160 => (x"de",x"4b",x"74",x"87"),
  1161 => (x"d8",x"ed",x"c2",x"93"),
  1162 => (x"49",x"a3",x"cb",x"83"),
  1163 => (x"84",x"c1",x"51",x"c0"),
  1164 => (x"cb",x"4a",x"6e",x"73"),
  1165 => (x"ef",x"f9",x"fe",x"49"),
  1166 => (x"48",x"66",x"c4",x"87"),
  1167 => (x"a6",x"c8",x"80",x"c1"),
  1168 => (x"03",x"ac",x"c7",x"58"),
  1169 => (x"6e",x"87",x"c5",x"c0"),
  1170 => (x"87",x"e0",x"fc",x"05"),
  1171 => (x"8e",x"f4",x"48",x"74"),
  1172 => (x"1e",x"87",x"fe",x"f5"),
  1173 => (x"4b",x"71",x"1e",x"73"),
  1174 => (x"c1",x"91",x"cb",x"49"),
  1175 => (x"c8",x"81",x"d4",x"e4"),
  1176 => (x"e4",x"c1",x"4a",x"a1"),
  1177 => (x"50",x"12",x"48",x"c0"),
  1178 => (x"c0",x"4a",x"a1",x"c9"),
  1179 => (x"12",x"48",x"dc",x"fa"),
  1180 => (x"c1",x"81",x"ca",x"50"),
  1181 => (x"11",x"48",x"c1",x"e4"),
  1182 => (x"c1",x"e4",x"c1",x"50"),
  1183 => (x"1e",x"49",x"bf",x"97"),
  1184 => (x"d3",x"f6",x"49",x"c0"),
  1185 => (x"ec",x"ec",x"c2",x"87"),
  1186 => (x"c1",x"78",x"de",x"48"),
  1187 => (x"87",x"d5",x"d6",x"49"),
  1188 => (x"87",x"c1",x"f5",x"26"),
  1189 => (x"49",x"4a",x"71",x"1e"),
  1190 => (x"e4",x"c1",x"91",x"cb"),
  1191 => (x"81",x"c8",x"81",x"d4"),
  1192 => (x"ec",x"c2",x"48",x"11"),
  1193 => (x"ed",x"c2",x"58",x"f0"),
  1194 => (x"78",x"c0",x"48",x"c4"),
  1195 => (x"f4",x"d5",x"49",x"c1"),
  1196 => (x"1e",x"4f",x"26",x"87"),
  1197 => (x"fe",x"c0",x"49",x"c0"),
  1198 => (x"4f",x"26",x"87",x"df"),
  1199 => (x"02",x"99",x"71",x"1e"),
  1200 => (x"e5",x"c1",x"87",x"d2"),
  1201 => (x"50",x"c0",x"48",x"e9"),
  1202 => (x"ca",x"c1",x"80",x"f7"),
  1203 => (x"e4",x"c1",x"40",x"d4"),
  1204 => (x"87",x"ce",x"78",x"cd"),
  1205 => (x"48",x"e5",x"e5",x"c1"),
  1206 => (x"78",x"c6",x"e4",x"c1"),
  1207 => (x"ca",x"c1",x"80",x"fc"),
  1208 => (x"4f",x"26",x"78",x"f3"),
  1209 => (x"5c",x"5b",x"5e",x"0e"),
  1210 => (x"4a",x"4c",x"71",x"0e"),
  1211 => (x"e4",x"c1",x"92",x"cb"),
  1212 => (x"a2",x"c8",x"82",x"d4"),
  1213 => (x"4b",x"a2",x"c9",x"49"),
  1214 => (x"1e",x"4b",x"6b",x"97"),
  1215 => (x"1e",x"49",x"69",x"97"),
  1216 => (x"49",x"12",x"82",x"ca"),
  1217 => (x"87",x"d8",x"e7",x"c0"),
  1218 => (x"d8",x"d4",x"49",x"c0"),
  1219 => (x"c0",x"49",x"74",x"87"),
  1220 => (x"f8",x"87",x"e1",x"fb"),
  1221 => (x"87",x"fb",x"f2",x"8e"),
  1222 => (x"71",x"1e",x"73",x"1e"),
  1223 => (x"c3",x"ff",x"49",x"4b"),
  1224 => (x"fe",x"49",x"73",x"87"),
  1225 => (x"ec",x"f2",x"87",x"fe"),
  1226 => (x"1e",x"73",x"1e",x"87"),
  1227 => (x"a3",x"c6",x"4b",x"71"),
  1228 => (x"87",x"db",x"02",x"4a"),
  1229 => (x"d6",x"02",x"8a",x"c1"),
  1230 => (x"c1",x"02",x"8a",x"87"),
  1231 => (x"02",x"8a",x"87",x"da"),
  1232 => (x"8a",x"87",x"fc",x"c0"),
  1233 => (x"87",x"e1",x"c0",x"02"),
  1234 => (x"87",x"cb",x"02",x"8a"),
  1235 => (x"c7",x"87",x"db",x"c1"),
  1236 => (x"87",x"c0",x"fd",x"49"),
  1237 => (x"c2",x"87",x"de",x"c1"),
  1238 => (x"02",x"bf",x"c4",x"ed"),
  1239 => (x"48",x"87",x"cb",x"c1"),
  1240 => (x"ed",x"c2",x"88",x"c1"),
  1241 => (x"c1",x"c1",x"58",x"c8"),
  1242 => (x"c8",x"ed",x"c2",x"87"),
  1243 => (x"f9",x"c0",x"02",x"bf"),
  1244 => (x"c4",x"ed",x"c2",x"87"),
  1245 => (x"80",x"c1",x"48",x"bf"),
  1246 => (x"58",x"c8",x"ed",x"c2"),
  1247 => (x"c2",x"87",x"eb",x"c0"),
  1248 => (x"49",x"bf",x"c4",x"ed"),
  1249 => (x"ed",x"c2",x"89",x"c6"),
  1250 => (x"b7",x"c0",x"59",x"c8"),
  1251 => (x"87",x"da",x"03",x"a9"),
  1252 => (x"48",x"c4",x"ed",x"c2"),
  1253 => (x"87",x"d2",x"78",x"c0"),
  1254 => (x"bf",x"c8",x"ed",x"c2"),
  1255 => (x"c2",x"87",x"cb",x"02"),
  1256 => (x"48",x"bf",x"c4",x"ed"),
  1257 => (x"ed",x"c2",x"80",x"c6"),
  1258 => (x"49",x"c0",x"58",x"c8"),
  1259 => (x"73",x"87",x"f6",x"d1"),
  1260 => (x"ff",x"f8",x"c0",x"49"),
  1261 => (x"87",x"dd",x"f0",x"87"),
  1262 => (x"5c",x"5b",x"5e",x"0e"),
  1263 => (x"d0",x"ff",x"0e",x"5d"),
  1264 => (x"59",x"a6",x"dc",x"86"),
  1265 => (x"c0",x"48",x"a6",x"c8"),
  1266 => (x"c1",x"80",x"c4",x"78"),
  1267 => (x"c4",x"78",x"66",x"c4"),
  1268 => (x"c4",x"78",x"c1",x"80"),
  1269 => (x"c2",x"78",x"c1",x"80"),
  1270 => (x"c1",x"48",x"c8",x"ed"),
  1271 => (x"ec",x"ec",x"c2",x"78"),
  1272 => (x"a8",x"de",x"48",x"bf"),
  1273 => (x"f4",x"87",x"cb",x"05"),
  1274 => (x"49",x"70",x"87",x"db"),
  1275 => (x"cf",x"59",x"a6",x"cc"),
  1276 => (x"e2",x"e3",x"87",x"f2"),
  1277 => (x"87",x"c4",x"e4",x"87"),
  1278 => (x"70",x"87",x"d1",x"e3"),
  1279 => (x"ac",x"fb",x"c0",x"4c"),
  1280 => (x"87",x"fb",x"c1",x"02"),
  1281 => (x"c1",x"05",x"66",x"d8"),
  1282 => (x"c0",x"c1",x"87",x"ed"),
  1283 => (x"82",x"c4",x"4a",x"66"),
  1284 => (x"1e",x"72",x"7e",x"6a"),
  1285 => (x"48",x"d9",x"e0",x"c1"),
  1286 => (x"c8",x"49",x"66",x"c4"),
  1287 => (x"41",x"20",x"4a",x"a1"),
  1288 => (x"f9",x"05",x"aa",x"71"),
  1289 => (x"26",x"51",x"10",x"87"),
  1290 => (x"66",x"c0",x"c1",x"4a"),
  1291 => (x"d3",x"c9",x"c1",x"48"),
  1292 => (x"c7",x"49",x"6a",x"78"),
  1293 => (x"c1",x"51",x"74",x"81"),
  1294 => (x"c8",x"49",x"66",x"c0"),
  1295 => (x"c1",x"51",x"c1",x"81"),
  1296 => (x"c9",x"49",x"66",x"c0"),
  1297 => (x"c1",x"51",x"c0",x"81"),
  1298 => (x"ca",x"49",x"66",x"c0"),
  1299 => (x"c1",x"51",x"c0",x"81"),
  1300 => (x"6a",x"1e",x"d8",x"1e"),
  1301 => (x"e2",x"81",x"c8",x"49"),
  1302 => (x"86",x"c8",x"87",x"f6"),
  1303 => (x"48",x"66",x"c4",x"c1"),
  1304 => (x"c7",x"01",x"a8",x"c0"),
  1305 => (x"48",x"a6",x"c8",x"87"),
  1306 => (x"87",x"ce",x"78",x"c1"),
  1307 => (x"48",x"66",x"c4",x"c1"),
  1308 => (x"a6",x"d0",x"88",x"c1"),
  1309 => (x"e2",x"87",x"c3",x"58"),
  1310 => (x"a6",x"d0",x"87",x"c2"),
  1311 => (x"74",x"78",x"c2",x"48"),
  1312 => (x"db",x"cd",x"02",x"9c"),
  1313 => (x"48",x"66",x"c8",x"87"),
  1314 => (x"a8",x"66",x"c8",x"c1"),
  1315 => (x"87",x"d0",x"cd",x"03"),
  1316 => (x"c0",x"48",x"a6",x"dc"),
  1317 => (x"c0",x"80",x"e8",x"78"),
  1318 => (x"87",x"f0",x"e0",x"78"),
  1319 => (x"d0",x"c1",x"4c",x"70"),
  1320 => (x"d9",x"c2",x"05",x"ac"),
  1321 => (x"7e",x"66",x"c4",x"87"),
  1322 => (x"70",x"87",x"d4",x"e3"),
  1323 => (x"59",x"a6",x"c8",x"49"),
  1324 => (x"70",x"87",x"d9",x"e0"),
  1325 => (x"ac",x"ec",x"c0",x"4c"),
  1326 => (x"87",x"ed",x"c1",x"05"),
  1327 => (x"cb",x"49",x"66",x"c8"),
  1328 => (x"66",x"c0",x"c1",x"91"),
  1329 => (x"4a",x"a1",x"c4",x"81"),
  1330 => (x"a1",x"c8",x"4d",x"6a"),
  1331 => (x"52",x"66",x"c4",x"4a"),
  1332 => (x"79",x"d4",x"ca",x"c1"),
  1333 => (x"87",x"f4",x"df",x"ff"),
  1334 => (x"02",x"9c",x"4c",x"70"),
  1335 => (x"fb",x"c0",x"87",x"d9"),
  1336 => (x"87",x"d3",x"02",x"ac"),
  1337 => (x"df",x"ff",x"55",x"74"),
  1338 => (x"4c",x"70",x"87",x"e2"),
  1339 => (x"87",x"c7",x"02",x"9c"),
  1340 => (x"05",x"ac",x"fb",x"c0"),
  1341 => (x"c0",x"87",x"ed",x"ff"),
  1342 => (x"c1",x"c2",x"55",x"e0"),
  1343 => (x"7d",x"97",x"c0",x"55"),
  1344 => (x"6e",x"49",x"66",x"d8"),
  1345 => (x"87",x"db",x"05",x"a9"),
  1346 => (x"cc",x"48",x"66",x"c8"),
  1347 => (x"ca",x"04",x"a8",x"66"),
  1348 => (x"48",x"66",x"c8",x"87"),
  1349 => (x"a6",x"cc",x"80",x"c1"),
  1350 => (x"cc",x"87",x"c8",x"58"),
  1351 => (x"88",x"c1",x"48",x"66"),
  1352 => (x"ff",x"58",x"a6",x"d0"),
  1353 => (x"70",x"87",x"e5",x"de"),
  1354 => (x"ac",x"d0",x"c1",x"4c"),
  1355 => (x"d4",x"87",x"c8",x"05"),
  1356 => (x"80",x"c1",x"48",x"66"),
  1357 => (x"c1",x"58",x"a6",x"d8"),
  1358 => (x"fd",x"02",x"ac",x"d0"),
  1359 => (x"e0",x"c0",x"87",x"e7"),
  1360 => (x"66",x"d8",x"48",x"a6"),
  1361 => (x"48",x"66",x"c4",x"78"),
  1362 => (x"a8",x"66",x"e0",x"c0"),
  1363 => (x"87",x"e2",x"c9",x"05"),
  1364 => (x"48",x"a6",x"e4",x"c0"),
  1365 => (x"80",x"c4",x"78",x"c0"),
  1366 => (x"48",x"74",x"78",x"c0"),
  1367 => (x"70",x"88",x"fb",x"c0"),
  1368 => (x"c8",x"02",x"6e",x"7e"),
  1369 => (x"48",x"6e",x"87",x"e5"),
  1370 => (x"7e",x"70",x"88",x"cb"),
  1371 => (x"cd",x"c1",x"02",x"6e"),
  1372 => (x"c9",x"48",x"6e",x"87"),
  1373 => (x"6e",x"7e",x"70",x"88"),
  1374 => (x"87",x"e9",x"c3",x"02"),
  1375 => (x"88",x"c4",x"48",x"6e"),
  1376 => (x"02",x"6e",x"7e",x"70"),
  1377 => (x"48",x"6e",x"87",x"ce"),
  1378 => (x"7e",x"70",x"88",x"c1"),
  1379 => (x"d4",x"c3",x"02",x"6e"),
  1380 => (x"87",x"f1",x"c7",x"87"),
  1381 => (x"c0",x"48",x"a6",x"dc"),
  1382 => (x"dc",x"ff",x"78",x"f0"),
  1383 => (x"4c",x"70",x"87",x"ee"),
  1384 => (x"02",x"ac",x"ec",x"c0"),
  1385 => (x"c0",x"87",x"c4",x"c0"),
  1386 => (x"c0",x"5c",x"a6",x"e0"),
  1387 => (x"cd",x"02",x"ac",x"ec"),
  1388 => (x"d7",x"dc",x"ff",x"87"),
  1389 => (x"c0",x"4c",x"70",x"87"),
  1390 => (x"ff",x"05",x"ac",x"ec"),
  1391 => (x"ec",x"c0",x"87",x"f3"),
  1392 => (x"c4",x"c0",x"02",x"ac"),
  1393 => (x"c3",x"dc",x"ff",x"87"),
  1394 => (x"ca",x"1e",x"c0",x"87"),
  1395 => (x"49",x"66",x"d0",x"1e"),
  1396 => (x"c8",x"c1",x"91",x"cb"),
  1397 => (x"80",x"71",x"48",x"66"),
  1398 => (x"c8",x"58",x"a6",x"cc"),
  1399 => (x"80",x"c4",x"48",x"66"),
  1400 => (x"cc",x"58",x"a6",x"d0"),
  1401 => (x"ff",x"49",x"bf",x"66"),
  1402 => (x"c1",x"87",x"e5",x"dc"),
  1403 => (x"d4",x"1e",x"de",x"1e"),
  1404 => (x"ff",x"49",x"bf",x"66"),
  1405 => (x"d0",x"87",x"d9",x"dc"),
  1406 => (x"c0",x"49",x"70",x"86"),
  1407 => (x"ec",x"c0",x"89",x"09"),
  1408 => (x"e8",x"c0",x"59",x"a6"),
  1409 => (x"a8",x"c0",x"48",x"66"),
  1410 => (x"87",x"ee",x"c0",x"06"),
  1411 => (x"48",x"66",x"e8",x"c0"),
  1412 => (x"c0",x"03",x"a8",x"dd"),
  1413 => (x"66",x"c4",x"87",x"e4"),
  1414 => (x"e8",x"c0",x"49",x"bf"),
  1415 => (x"e0",x"c0",x"81",x"66"),
  1416 => (x"66",x"e8",x"c0",x"51"),
  1417 => (x"c4",x"81",x"c1",x"49"),
  1418 => (x"c2",x"81",x"bf",x"66"),
  1419 => (x"e8",x"c0",x"51",x"c1"),
  1420 => (x"81",x"c2",x"49",x"66"),
  1421 => (x"81",x"bf",x"66",x"c4"),
  1422 => (x"48",x"6e",x"51",x"c0"),
  1423 => (x"78",x"d3",x"c9",x"c1"),
  1424 => (x"81",x"c8",x"49",x"6e"),
  1425 => (x"6e",x"51",x"66",x"d0"),
  1426 => (x"d4",x"81",x"c9",x"49"),
  1427 => (x"49",x"6e",x"51",x"66"),
  1428 => (x"66",x"dc",x"81",x"ca"),
  1429 => (x"48",x"66",x"d0",x"51"),
  1430 => (x"a6",x"d4",x"80",x"c1"),
  1431 => (x"80",x"d8",x"48",x"58"),
  1432 => (x"e6",x"c4",x"78",x"c1"),
  1433 => (x"d6",x"dc",x"ff",x"87"),
  1434 => (x"c0",x"49",x"70",x"87"),
  1435 => (x"ff",x"59",x"a6",x"ec"),
  1436 => (x"70",x"87",x"cc",x"dc"),
  1437 => (x"a6",x"e0",x"c0",x"49"),
  1438 => (x"48",x"66",x"dc",x"59"),
  1439 => (x"05",x"a8",x"ec",x"c0"),
  1440 => (x"dc",x"87",x"ca",x"c0"),
  1441 => (x"e8",x"c0",x"48",x"a6"),
  1442 => (x"c4",x"c0",x"78",x"66"),
  1443 => (x"fb",x"d8",x"ff",x"87"),
  1444 => (x"49",x"66",x"c8",x"87"),
  1445 => (x"c0",x"c1",x"91",x"cb"),
  1446 => (x"80",x"71",x"48",x"66"),
  1447 => (x"49",x"6e",x"7e",x"70"),
  1448 => (x"4a",x"6e",x"81",x"c8"),
  1449 => (x"e8",x"c0",x"82",x"ca"),
  1450 => (x"66",x"dc",x"52",x"66"),
  1451 => (x"c0",x"82",x"c1",x"4a"),
  1452 => (x"c1",x"8a",x"66",x"e8"),
  1453 => (x"70",x"30",x"72",x"48"),
  1454 => (x"72",x"8a",x"c1",x"4a"),
  1455 => (x"69",x"97",x"79",x"97"),
  1456 => (x"ec",x"c0",x"1e",x"49"),
  1457 => (x"d9",x"d7",x"49",x"66"),
  1458 => (x"c0",x"86",x"c4",x"87"),
  1459 => (x"6e",x"58",x"a6",x"f0"),
  1460 => (x"69",x"81",x"c4",x"49"),
  1461 => (x"66",x"e0",x"c0",x"4d"),
  1462 => (x"a8",x"66",x"c4",x"48"),
  1463 => (x"87",x"c8",x"c0",x"02"),
  1464 => (x"c0",x"48",x"a6",x"c4"),
  1465 => (x"87",x"c5",x"c0",x"78"),
  1466 => (x"c1",x"48",x"a6",x"c4"),
  1467 => (x"1e",x"66",x"c4",x"78"),
  1468 => (x"75",x"1e",x"e0",x"c0"),
  1469 => (x"d7",x"d8",x"ff",x"49"),
  1470 => (x"70",x"86",x"c8",x"87"),
  1471 => (x"ac",x"b7",x"c0",x"4c"),
  1472 => (x"87",x"d4",x"c1",x"06"),
  1473 => (x"e0",x"c0",x"85",x"74"),
  1474 => (x"75",x"89",x"74",x"49"),
  1475 => (x"e2",x"e0",x"c1",x"4b"),
  1476 => (x"e6",x"fe",x"71",x"4a"),
  1477 => (x"85",x"c2",x"87",x"d2"),
  1478 => (x"48",x"66",x"e4",x"c0"),
  1479 => (x"e8",x"c0",x"80",x"c1"),
  1480 => (x"ec",x"c0",x"58",x"a6"),
  1481 => (x"81",x"c1",x"49",x"66"),
  1482 => (x"c0",x"02",x"a9",x"70"),
  1483 => (x"a6",x"c4",x"87",x"c8"),
  1484 => (x"c0",x"78",x"c0",x"48"),
  1485 => (x"a6",x"c4",x"87",x"c5"),
  1486 => (x"c4",x"78",x"c1",x"48"),
  1487 => (x"a4",x"c2",x"1e",x"66"),
  1488 => (x"48",x"e0",x"c0",x"49"),
  1489 => (x"49",x"70",x"88",x"71"),
  1490 => (x"ff",x"49",x"75",x"1e"),
  1491 => (x"c8",x"87",x"c1",x"d7"),
  1492 => (x"a8",x"b7",x"c0",x"86"),
  1493 => (x"87",x"c0",x"ff",x"01"),
  1494 => (x"02",x"66",x"e4",x"c0"),
  1495 => (x"6e",x"87",x"d1",x"c0"),
  1496 => (x"c0",x"81",x"c9",x"49"),
  1497 => (x"6e",x"51",x"66",x"e4"),
  1498 => (x"e4",x"cb",x"c1",x"48"),
  1499 => (x"87",x"cc",x"c0",x"78"),
  1500 => (x"81",x"c9",x"49",x"6e"),
  1501 => (x"48",x"6e",x"51",x"c2"),
  1502 => (x"78",x"d8",x"cc",x"c1"),
  1503 => (x"48",x"a6",x"e8",x"c0"),
  1504 => (x"c6",x"c0",x"78",x"c1"),
  1505 => (x"f3",x"d5",x"ff",x"87"),
  1506 => (x"c0",x"4c",x"70",x"87"),
  1507 => (x"c0",x"02",x"66",x"e8"),
  1508 => (x"66",x"c8",x"87",x"f5"),
  1509 => (x"a8",x"66",x"cc",x"48"),
  1510 => (x"87",x"cb",x"c0",x"04"),
  1511 => (x"c1",x"48",x"66",x"c8"),
  1512 => (x"58",x"a6",x"cc",x"80"),
  1513 => (x"cc",x"87",x"e0",x"c0"),
  1514 => (x"88",x"c1",x"48",x"66"),
  1515 => (x"c0",x"58",x"a6",x"d0"),
  1516 => (x"c6",x"c1",x"87",x"d5"),
  1517 => (x"c8",x"c0",x"05",x"ac"),
  1518 => (x"48",x"66",x"d0",x"87"),
  1519 => (x"a6",x"d4",x"80",x"c1"),
  1520 => (x"f7",x"d4",x"ff",x"58"),
  1521 => (x"d4",x"4c",x"70",x"87"),
  1522 => (x"80",x"c1",x"48",x"66"),
  1523 => (x"74",x"58",x"a6",x"d8"),
  1524 => (x"cb",x"c0",x"02",x"9c"),
  1525 => (x"48",x"66",x"c8",x"87"),
  1526 => (x"a8",x"66",x"c8",x"c1"),
  1527 => (x"87",x"f0",x"f2",x"04"),
  1528 => (x"87",x"cf",x"d4",x"ff"),
  1529 => (x"c7",x"48",x"66",x"c8"),
  1530 => (x"e5",x"c0",x"03",x"a8"),
  1531 => (x"c8",x"ed",x"c2",x"87"),
  1532 => (x"c8",x"78",x"c0",x"48"),
  1533 => (x"91",x"cb",x"49",x"66"),
  1534 => (x"81",x"66",x"c0",x"c1"),
  1535 => (x"6a",x"4a",x"a1",x"c4"),
  1536 => (x"79",x"52",x"c0",x"4a"),
  1537 => (x"c1",x"48",x"66",x"c8"),
  1538 => (x"58",x"a6",x"cc",x"80"),
  1539 => (x"ff",x"04",x"a8",x"c7"),
  1540 => (x"d0",x"ff",x"87",x"db"),
  1541 => (x"f8",x"de",x"ff",x"8e"),
  1542 => (x"61",x"6f",x"4c",x"87"),
  1543 => (x"2e",x"2a",x"20",x"64"),
  1544 => (x"20",x"3a",x"00",x"20"),
  1545 => (x"1e",x"73",x"1e",x"00"),
  1546 => (x"02",x"9b",x"4b",x"71"),
  1547 => (x"ed",x"c2",x"87",x"c6"),
  1548 => (x"78",x"c0",x"48",x"c4"),
  1549 => (x"ed",x"c2",x"1e",x"c7"),
  1550 => (x"1e",x"49",x"bf",x"c4"),
  1551 => (x"1e",x"d4",x"e4",x"c1"),
  1552 => (x"bf",x"ec",x"ec",x"c2"),
  1553 => (x"87",x"f0",x"ed",x"49"),
  1554 => (x"ec",x"c2",x"86",x"cc"),
  1555 => (x"e9",x"49",x"bf",x"ec"),
  1556 => (x"9b",x"73",x"87",x"ea"),
  1557 => (x"c1",x"87",x"c8",x"02"),
  1558 => (x"c0",x"49",x"d4",x"e4"),
  1559 => (x"ff",x"87",x"e7",x"e7"),
  1560 => (x"1e",x"87",x"f2",x"dd"),
  1561 => (x"48",x"c0",x"e4",x"c1"),
  1562 => (x"e5",x"c1",x"50",x"c0"),
  1563 => (x"ff",x"49",x"bf",x"f7"),
  1564 => (x"c0",x"87",x"ea",x"d8"),
  1565 => (x"1e",x"4f",x"26",x"48"),
  1566 => (x"c1",x"87",x"e3",x"c7"),
  1567 => (x"87",x"e5",x"fe",x"49"),
  1568 => (x"87",x"cc",x"e9",x"fe"),
  1569 => (x"cd",x"02",x"98",x"70"),
  1570 => (x"c7",x"f2",x"fe",x"87"),
  1571 => (x"02",x"98",x"70",x"87"),
  1572 => (x"4a",x"c1",x"87",x"c4"),
  1573 => (x"4a",x"c0",x"87",x"c2"),
  1574 => (x"ce",x"05",x"9a",x"72"),
  1575 => (x"c1",x"1e",x"c0",x"87"),
  1576 => (x"c0",x"49",x"c7",x"e3"),
  1577 => (x"c4",x"87",x"f7",x"f2"),
  1578 => (x"c0",x"87",x"fe",x"86"),
  1579 => (x"d2",x"e3",x"c1",x"1e"),
  1580 => (x"e9",x"f2",x"c0",x"49"),
  1581 => (x"fe",x"1e",x"c0",x"87"),
  1582 => (x"49",x"70",x"87",x"e9"),
  1583 => (x"87",x"de",x"f2",x"c0"),
  1584 => (x"f8",x"87",x"da",x"c3"),
  1585 => (x"53",x"4f",x"26",x"8e"),
  1586 => (x"61",x"66",x"20",x"44"),
  1587 => (x"64",x"65",x"6c",x"69"),
  1588 => (x"6f",x"42",x"00",x"2e"),
  1589 => (x"6e",x"69",x"74",x"6f"),
  1590 => (x"2e",x"2e",x"2e",x"67"),
  1591 => (x"ea",x"c0",x"1e",x"00"),
  1592 => (x"f5",x"c0",x"87",x"c0"),
  1593 => (x"87",x"f6",x"87",x"ee"),
  1594 => (x"c2",x"1e",x"4f",x"26"),
  1595 => (x"c0",x"48",x"c4",x"ed"),
  1596 => (x"ec",x"ec",x"c2",x"78"),
  1597 => (x"fd",x"78",x"c0",x"48"),
  1598 => (x"87",x"e1",x"87",x"fd"),
  1599 => (x"4f",x"26",x"48",x"c0"),
  1600 => (x"00",x"01",x"00",x"00"),
  1601 => (x"20",x"80",x"00",x"00"),
  1602 => (x"74",x"69",x"78",x"45"),
  1603 => (x"42",x"20",x"80",x"00"),
  1604 => (x"00",x"6b",x"63",x"61"),
  1605 => (x"00",x"00",x"12",x"94"),
  1606 => (x"00",x"00",x"2b",x"58"),
  1607 => (x"94",x"00",x"00",x"00"),
  1608 => (x"76",x"00",x"00",x"12"),
  1609 => (x"00",x"00",x"00",x"2b"),
  1610 => (x"12",x"94",x"00",x"00"),
  1611 => (x"2b",x"94",x"00",x"00"),
  1612 => (x"00",x"00",x"00",x"00"),
  1613 => (x"00",x"12",x"94",x"00"),
  1614 => (x"00",x"2b",x"b2",x"00"),
  1615 => (x"00",x"00",x"00",x"00"),
  1616 => (x"00",x"00",x"12",x"94"),
  1617 => (x"00",x"00",x"2b",x"d0"),
  1618 => (x"94",x"00",x"00",x"00"),
  1619 => (x"ee",x"00",x"00",x"12"),
  1620 => (x"00",x"00",x"00",x"2b"),
  1621 => (x"12",x"94",x"00",x"00"),
  1622 => (x"2c",x"0c",x"00",x"00"),
  1623 => (x"00",x"00",x"00",x"00"),
  1624 => (x"00",x"12",x"94",x"00"),
  1625 => (x"00",x"00",x"00",x"00"),
  1626 => (x"00",x"00",x"00",x"00"),
  1627 => (x"00",x"00",x"13",x"29"),
  1628 => (x"00",x"00",x"00",x"00"),
  1629 => (x"7b",x"00",x"00",x"00"),
  1630 => (x"43",x"00",x"00",x"19"),
  1631 => (x"20",x"20",x"34",x"36"),
  1632 => (x"52",x"20",x"20",x"20"),
  1633 => (x"1e",x"00",x"4d",x"4f"),
  1634 => (x"c0",x"48",x"f0",x"fe"),
  1635 => (x"79",x"09",x"cd",x"78"),
  1636 => (x"1e",x"4f",x"26",x"09"),
  1637 => (x"bf",x"f0",x"fe",x"1e"),
  1638 => (x"26",x"26",x"48",x"7e"),
  1639 => (x"f0",x"fe",x"1e",x"4f"),
  1640 => (x"26",x"78",x"c1",x"48"),
  1641 => (x"f0",x"fe",x"1e",x"4f"),
  1642 => (x"26",x"78",x"c0",x"48"),
  1643 => (x"4a",x"71",x"1e",x"4f"),
  1644 => (x"26",x"52",x"52",x"c0"),
  1645 => (x"5b",x"5e",x"0e",x"4f"),
  1646 => (x"f4",x"0e",x"5d",x"5c"),
  1647 => (x"97",x"4d",x"71",x"86"),
  1648 => (x"a5",x"c1",x"7e",x"6d"),
  1649 => (x"48",x"6c",x"97",x"4c"),
  1650 => (x"6e",x"58",x"a6",x"c8"),
  1651 => (x"a8",x"66",x"c4",x"48"),
  1652 => (x"ff",x"87",x"c5",x"05"),
  1653 => (x"87",x"e6",x"c0",x"48"),
  1654 => (x"c2",x"87",x"ca",x"ff"),
  1655 => (x"6c",x"97",x"49",x"a5"),
  1656 => (x"4b",x"a3",x"71",x"4b"),
  1657 => (x"97",x"4b",x"6b",x"97"),
  1658 => (x"48",x"6e",x"7e",x"6c"),
  1659 => (x"a6",x"c8",x"80",x"c1"),
  1660 => (x"cc",x"98",x"c7",x"58"),
  1661 => (x"97",x"70",x"58",x"a6"),
  1662 => (x"87",x"e1",x"fe",x"7c"),
  1663 => (x"8e",x"f4",x"48",x"73"),
  1664 => (x"4c",x"26",x"4d",x"26"),
  1665 => (x"4f",x"26",x"4b",x"26"),
  1666 => (x"5c",x"5b",x"5e",x"0e"),
  1667 => (x"71",x"86",x"f4",x"0e"),
  1668 => (x"4a",x"66",x"d8",x"4c"),
  1669 => (x"c2",x"9a",x"ff",x"c3"),
  1670 => (x"6c",x"97",x"4b",x"a4"),
  1671 => (x"49",x"a1",x"73",x"49"),
  1672 => (x"6c",x"97",x"51",x"72"),
  1673 => (x"c1",x"48",x"6e",x"7e"),
  1674 => (x"58",x"a6",x"c8",x"80"),
  1675 => (x"a6",x"cc",x"98",x"c7"),
  1676 => (x"f4",x"54",x"70",x"58"),
  1677 => (x"87",x"ca",x"ff",x"8e"),
  1678 => (x"e8",x"fd",x"1e",x"1e"),
  1679 => (x"4a",x"bf",x"e0",x"87"),
  1680 => (x"c0",x"e0",x"c0",x"49"),
  1681 => (x"87",x"cb",x"02",x"99"),
  1682 => (x"f0",x"c2",x"1e",x"72"),
  1683 => (x"f7",x"fe",x"49",x"ea"),
  1684 => (x"fc",x"86",x"c4",x"87"),
  1685 => (x"7e",x"70",x"87",x"fd"),
  1686 => (x"26",x"87",x"c2",x"fd"),
  1687 => (x"c2",x"1e",x"4f",x"26"),
  1688 => (x"fd",x"49",x"ea",x"f0"),
  1689 => (x"e8",x"c1",x"87",x"c7"),
  1690 => (x"da",x"fc",x"49",x"f8"),
  1691 => (x"87",x"c7",x"c4",x"87"),
  1692 => (x"ff",x"1e",x"4f",x"26"),
  1693 => (x"e1",x"c8",x"48",x"d0"),
  1694 => (x"48",x"d4",x"ff",x"78"),
  1695 => (x"66",x"c4",x"78",x"c5"),
  1696 => (x"c3",x"87",x"c3",x"02"),
  1697 => (x"66",x"c8",x"78",x"e0"),
  1698 => (x"ff",x"87",x"c6",x"02"),
  1699 => (x"f0",x"c3",x"48",x"d4"),
  1700 => (x"48",x"d4",x"ff",x"78"),
  1701 => (x"d0",x"ff",x"78",x"71"),
  1702 => (x"78",x"e1",x"c8",x"48"),
  1703 => (x"26",x"78",x"e0",x"c0"),
  1704 => (x"5b",x"5e",x"0e",x"4f"),
  1705 => (x"4c",x"71",x"0e",x"5c"),
  1706 => (x"49",x"ea",x"f0",x"c2"),
  1707 => (x"70",x"87",x"c6",x"fc"),
  1708 => (x"aa",x"b7",x"c0",x"4a"),
  1709 => (x"87",x"e2",x"c2",x"04"),
  1710 => (x"05",x"aa",x"f0",x"c3"),
  1711 => (x"ed",x"c1",x"87",x"c9"),
  1712 => (x"78",x"c1",x"48",x"e6"),
  1713 => (x"c3",x"87",x"c3",x"c2"),
  1714 => (x"c9",x"05",x"aa",x"e0"),
  1715 => (x"ea",x"ed",x"c1",x"87"),
  1716 => (x"c1",x"78",x"c1",x"48"),
  1717 => (x"ed",x"c1",x"87",x"f4"),
  1718 => (x"c6",x"02",x"bf",x"ea"),
  1719 => (x"a2",x"c0",x"c2",x"87"),
  1720 => (x"72",x"87",x"c2",x"4b"),
  1721 => (x"05",x"9c",x"74",x"4b"),
  1722 => (x"ed",x"c1",x"87",x"d1"),
  1723 => (x"c1",x"1e",x"bf",x"e6"),
  1724 => (x"1e",x"bf",x"ea",x"ed"),
  1725 => (x"f9",x"fd",x"49",x"72"),
  1726 => (x"c1",x"86",x"c8",x"87"),
  1727 => (x"02",x"bf",x"e6",x"ed"),
  1728 => (x"73",x"87",x"e0",x"c0"),
  1729 => (x"29",x"b7",x"c4",x"49"),
  1730 => (x"c6",x"ef",x"c1",x"91"),
  1731 => (x"cf",x"4a",x"73",x"81"),
  1732 => (x"c1",x"92",x"c2",x"9a"),
  1733 => (x"70",x"30",x"72",x"48"),
  1734 => (x"72",x"ba",x"ff",x"4a"),
  1735 => (x"70",x"98",x"69",x"48"),
  1736 => (x"73",x"87",x"db",x"79"),
  1737 => (x"29",x"b7",x"c4",x"49"),
  1738 => (x"c6",x"ef",x"c1",x"91"),
  1739 => (x"cf",x"4a",x"73",x"81"),
  1740 => (x"c3",x"92",x"c2",x"9a"),
  1741 => (x"70",x"30",x"72",x"48"),
  1742 => (x"b0",x"69",x"48",x"4a"),
  1743 => (x"ed",x"c1",x"79",x"70"),
  1744 => (x"78",x"c0",x"48",x"ea"),
  1745 => (x"48",x"e6",x"ed",x"c1"),
  1746 => (x"f0",x"c2",x"78",x"c0"),
  1747 => (x"e4",x"f9",x"49",x"ea"),
  1748 => (x"c0",x"4a",x"70",x"87"),
  1749 => (x"fd",x"03",x"aa",x"b7"),
  1750 => (x"48",x"c0",x"87",x"de"),
  1751 => (x"4d",x"26",x"87",x"c2"),
  1752 => (x"4b",x"26",x"4c",x"26"),
  1753 => (x"00",x"00",x"4f",x"26"),
  1754 => (x"00",x"00",x"00",x"00"),
  1755 => (x"71",x"1e",x"00",x"00"),
  1756 => (x"ec",x"fc",x"49",x"4a"),
  1757 => (x"1e",x"4f",x"26",x"87"),
  1758 => (x"49",x"72",x"4a",x"c0"),
  1759 => (x"ef",x"c1",x"91",x"c4"),
  1760 => (x"79",x"c0",x"81",x"c6"),
  1761 => (x"b7",x"d0",x"82",x"c1"),
  1762 => (x"87",x"ee",x"04",x"aa"),
  1763 => (x"5e",x"0e",x"4f",x"26"),
  1764 => (x"0e",x"5d",x"5c",x"5b"),
  1765 => (x"cc",x"f8",x"4d",x"71"),
  1766 => (x"c4",x"4a",x"75",x"87"),
  1767 => (x"c1",x"92",x"2a",x"b7"),
  1768 => (x"75",x"82",x"c6",x"ef"),
  1769 => (x"c2",x"9c",x"cf",x"4c"),
  1770 => (x"4b",x"49",x"6a",x"94"),
  1771 => (x"9b",x"c3",x"2b",x"74"),
  1772 => (x"30",x"74",x"48",x"c2"),
  1773 => (x"bc",x"ff",x"4c",x"70"),
  1774 => (x"98",x"71",x"48",x"74"),
  1775 => (x"dc",x"f7",x"7a",x"70"),
  1776 => (x"fe",x"48",x"73",x"87"),
  1777 => (x"00",x"00",x"87",x"d8"),
  1778 => (x"00",x"00",x"00",x"00"),
  1779 => (x"00",x"00",x"00",x"00"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"00",x"00",x"00",x"00"),
  1784 => (x"00",x"00",x"00",x"00"),
  1785 => (x"00",x"00",x"00",x"00"),
  1786 => (x"00",x"00",x"00",x"00"),
  1787 => (x"00",x"00",x"00",x"00"),
  1788 => (x"00",x"00",x"00",x"00"),
  1789 => (x"00",x"00",x"00",x"00"),
  1790 => (x"00",x"00",x"00",x"00"),
  1791 => (x"00",x"00",x"00",x"00"),
  1792 => (x"00",x"00",x"00",x"00"),
  1793 => (x"ff",x"1e",x"00",x"00"),
  1794 => (x"e1",x"c8",x"48",x"d0"),
  1795 => (x"ff",x"48",x"71",x"78"),
  1796 => (x"26",x"78",x"08",x"d4"),
  1797 => (x"d0",x"ff",x"1e",x"4f"),
  1798 => (x"78",x"e1",x"c8",x"48"),
  1799 => (x"d4",x"ff",x"48",x"71"),
  1800 => (x"66",x"c4",x"78",x"08"),
  1801 => (x"08",x"d4",x"ff",x"48"),
  1802 => (x"1e",x"4f",x"26",x"78"),
  1803 => (x"66",x"c4",x"4a",x"71"),
  1804 => (x"49",x"72",x"1e",x"49"),
  1805 => (x"ff",x"87",x"de",x"ff"),
  1806 => (x"e0",x"c0",x"48",x"d0"),
  1807 => (x"4f",x"26",x"26",x"78"),
  1808 => (x"71",x"1e",x"73",x"1e"),
  1809 => (x"49",x"66",x"c8",x"4b"),
  1810 => (x"c1",x"4a",x"73",x"1e"),
  1811 => (x"ff",x"49",x"a2",x"e0"),
  1812 => (x"c4",x"26",x"87",x"d9"),
  1813 => (x"26",x"4d",x"26",x"87"),
  1814 => (x"26",x"4b",x"26",x"4c"),
  1815 => (x"d4",x"ff",x"1e",x"4f"),
  1816 => (x"7a",x"ff",x"c3",x"4a"),
  1817 => (x"c0",x"48",x"d0",x"ff"),
  1818 => (x"7a",x"de",x"78",x"e1"),
  1819 => (x"bf",x"f4",x"f0",x"c2"),
  1820 => (x"c8",x"48",x"49",x"7a"),
  1821 => (x"71",x"7a",x"70",x"28"),
  1822 => (x"70",x"28",x"d0",x"48"),
  1823 => (x"d8",x"48",x"71",x"7a"),
  1824 => (x"c2",x"7a",x"70",x"28"),
  1825 => (x"7a",x"bf",x"f8",x"f0"),
  1826 => (x"28",x"c8",x"48",x"49"),
  1827 => (x"48",x"71",x"7a",x"70"),
  1828 => (x"7a",x"70",x"28",x"d0"),
  1829 => (x"28",x"d8",x"48",x"71"),
  1830 => (x"d0",x"ff",x"7a",x"70"),
  1831 => (x"78",x"e0",x"c0",x"48"),
  1832 => (x"73",x"1e",x"4f",x"26"),
  1833 => (x"c2",x"4a",x"71",x"1e"),
  1834 => (x"4b",x"bf",x"f4",x"f0"),
  1835 => (x"e0",x"c0",x"2b",x"72"),
  1836 => (x"87",x"ce",x"04",x"aa"),
  1837 => (x"e0",x"c0",x"49",x"72"),
  1838 => (x"f8",x"f0",x"c2",x"89"),
  1839 => (x"2b",x"71",x"4b",x"bf"),
  1840 => (x"e0",x"c0",x"87",x"cf"),
  1841 => (x"c2",x"89",x"72",x"49"),
  1842 => (x"48",x"bf",x"f8",x"f0"),
  1843 => (x"49",x"70",x"30",x"71"),
  1844 => (x"9b",x"66",x"c8",x"b3"),
  1845 => (x"87",x"c4",x"48",x"73"),
  1846 => (x"4c",x"26",x"4d",x"26"),
  1847 => (x"4f",x"26",x"4b",x"26"),
  1848 => (x"5c",x"5b",x"5e",x"0e"),
  1849 => (x"86",x"ec",x"0e",x"5d"),
  1850 => (x"f0",x"c2",x"4b",x"71"),
  1851 => (x"4c",x"7e",x"bf",x"f4"),
  1852 => (x"e0",x"c0",x"2c",x"73"),
  1853 => (x"e0",x"c0",x"04",x"ab"),
  1854 => (x"48",x"a6",x"c4",x"87"),
  1855 => (x"49",x"73",x"78",x"c0"),
  1856 => (x"71",x"89",x"e0",x"c0"),
  1857 => (x"66",x"e4",x"c0",x"4a"),
  1858 => (x"cc",x"30",x"72",x"48"),
  1859 => (x"f0",x"c2",x"58",x"a6"),
  1860 => (x"4c",x"4d",x"bf",x"f8"),
  1861 => (x"e4",x"c0",x"2c",x"71"),
  1862 => (x"c0",x"49",x"73",x"87"),
  1863 => (x"71",x"48",x"66",x"e4"),
  1864 => (x"58",x"a6",x"c8",x"30"),
  1865 => (x"73",x"49",x"e0",x"c0"),
  1866 => (x"66",x"e4",x"c0",x"89"),
  1867 => (x"cc",x"28",x"71",x"48"),
  1868 => (x"f0",x"c2",x"58",x"a6"),
  1869 => (x"48",x"4d",x"bf",x"f8"),
  1870 => (x"49",x"70",x"30",x"71"),
  1871 => (x"66",x"e4",x"c0",x"b4"),
  1872 => (x"c0",x"84",x"c1",x"9c"),
  1873 => (x"04",x"ac",x"66",x"e8"),
  1874 => (x"4c",x"c0",x"87",x"c2"),
  1875 => (x"04",x"ab",x"e0",x"c0"),
  1876 => (x"a6",x"cc",x"87",x"d3"),
  1877 => (x"73",x"78",x"c0",x"48"),
  1878 => (x"89",x"e0",x"c0",x"49"),
  1879 => (x"30",x"71",x"48",x"74"),
  1880 => (x"d5",x"58",x"a6",x"d4"),
  1881 => (x"74",x"49",x"73",x"87"),
  1882 => (x"d0",x"30",x"71",x"48"),
  1883 => (x"e0",x"c0",x"58",x"a6"),
  1884 => (x"74",x"89",x"73",x"49"),
  1885 => (x"d4",x"28",x"71",x"48"),
  1886 => (x"66",x"c4",x"58",x"a6"),
  1887 => (x"6e",x"ba",x"ff",x"4a"),
  1888 => (x"49",x"66",x"c8",x"9a"),
  1889 => (x"99",x"75",x"b9",x"ff"),
  1890 => (x"66",x"cc",x"48",x"72"),
  1891 => (x"f8",x"f0",x"c2",x"b0"),
  1892 => (x"d0",x"48",x"71",x"58"),
  1893 => (x"f0",x"c2",x"b0",x"66"),
  1894 => (x"c0",x"fb",x"58",x"fc"),
  1895 => (x"fc",x"8e",x"ec",x"87"),
  1896 => (x"ff",x"1e",x"87",x"f6"),
  1897 => (x"c9",x"c8",x"48",x"d0"),
  1898 => (x"ff",x"48",x"71",x"78"),
  1899 => (x"26",x"78",x"08",x"d4"),
  1900 => (x"4a",x"71",x"1e",x"4f"),
  1901 => (x"ff",x"87",x"eb",x"49"),
  1902 => (x"78",x"c8",x"48",x"d0"),
  1903 => (x"73",x"1e",x"4f",x"26"),
  1904 => (x"c2",x"4b",x"71",x"1e"),
  1905 => (x"02",x"bf",x"c8",x"f1"),
  1906 => (x"eb",x"c2",x"87",x"c3"),
  1907 => (x"48",x"d0",x"ff",x"87"),
  1908 => (x"73",x"78",x"c9",x"c8"),
  1909 => (x"b1",x"e0",x"c0",x"49"),
  1910 => (x"71",x"48",x"d4",x"ff"),
  1911 => (x"fc",x"f0",x"c2",x"78"),
  1912 => (x"c8",x"78",x"c0",x"48"),
  1913 => (x"87",x"c5",x"02",x"66"),
  1914 => (x"c2",x"49",x"ff",x"c3"),
  1915 => (x"c2",x"49",x"c0",x"87"),
  1916 => (x"cc",x"59",x"c4",x"f1"),
  1917 => (x"87",x"c6",x"02",x"66"),
  1918 => (x"4a",x"d5",x"d5",x"c5"),
  1919 => (x"ff",x"cf",x"87",x"c4"),
  1920 => (x"f1",x"c2",x"4a",x"ff"),
  1921 => (x"f1",x"c2",x"5a",x"c8"),
  1922 => (x"78",x"c1",x"48",x"c8"),
  1923 => (x"4d",x"26",x"87",x"c4"),
  1924 => (x"4b",x"26",x"4c",x"26"),
  1925 => (x"5e",x"0e",x"4f",x"26"),
  1926 => (x"0e",x"5d",x"5c",x"5b"),
  1927 => (x"f1",x"c2",x"4a",x"71"),
  1928 => (x"72",x"4c",x"bf",x"c4"),
  1929 => (x"87",x"cb",x"02",x"9a"),
  1930 => (x"c1",x"91",x"c8",x"49"),
  1931 => (x"71",x"4b",x"f4",x"f6"),
  1932 => (x"c1",x"87",x"c4",x"83"),
  1933 => (x"c0",x"4b",x"f4",x"fa"),
  1934 => (x"74",x"49",x"13",x"4d"),
  1935 => (x"c0",x"f1",x"c2",x"99"),
  1936 => (x"d4",x"ff",x"b9",x"bf"),
  1937 => (x"c1",x"78",x"71",x"48"),
  1938 => (x"c8",x"85",x"2c",x"b7"),
  1939 => (x"e8",x"04",x"ad",x"b7"),
  1940 => (x"fc",x"f0",x"c2",x"87"),
  1941 => (x"80",x"c8",x"48",x"bf"),
  1942 => (x"58",x"c0",x"f1",x"c2"),
  1943 => (x"1e",x"87",x"ef",x"fe"),
  1944 => (x"4b",x"71",x"1e",x"73"),
  1945 => (x"02",x"9a",x"4a",x"13"),
  1946 => (x"49",x"72",x"87",x"cb"),
  1947 => (x"13",x"87",x"e7",x"fe"),
  1948 => (x"f5",x"05",x"9a",x"4a"),
  1949 => (x"87",x"da",x"fe",x"87"),
  1950 => (x"fc",x"f0",x"c2",x"1e"),
  1951 => (x"f0",x"c2",x"49",x"bf"),
  1952 => (x"a1",x"c1",x"48",x"fc"),
  1953 => (x"b7",x"c0",x"c4",x"78"),
  1954 => (x"87",x"db",x"03",x"a9"),
  1955 => (x"c2",x"48",x"d4",x"ff"),
  1956 => (x"78",x"bf",x"c0",x"f1"),
  1957 => (x"bf",x"fc",x"f0",x"c2"),
  1958 => (x"fc",x"f0",x"c2",x"49"),
  1959 => (x"78",x"a1",x"c1",x"48"),
  1960 => (x"a9",x"b7",x"c0",x"c4"),
  1961 => (x"ff",x"87",x"e5",x"04"),
  1962 => (x"78",x"c8",x"48",x"d0"),
  1963 => (x"48",x"c8",x"f1",x"c2"),
  1964 => (x"4f",x"26",x"78",x"c0"),
  1965 => (x"00",x"00",x"00",x"00"),
  1966 => (x"00",x"00",x"00",x"00"),
  1967 => (x"5f",x"00",x"00",x"00"),
  1968 => (x"00",x"00",x"00",x"5f"),
  1969 => (x"00",x"03",x"03",x"00"),
  1970 => (x"00",x"00",x"03",x"03"),
  1971 => (x"14",x"7f",x"7f",x"14"),
  1972 => (x"00",x"14",x"7f",x"7f"),
  1973 => (x"6b",x"2e",x"24",x"00"),
  1974 => (x"00",x"12",x"3a",x"6b"),
  1975 => (x"18",x"36",x"6a",x"4c"),
  1976 => (x"00",x"32",x"56",x"6c"),
  1977 => (x"59",x"4f",x"7e",x"30"),
  1978 => (x"40",x"68",x"3a",x"77"),
  1979 => (x"07",x"04",x"00",x"00"),
  1980 => (x"00",x"00",x"00",x"03"),
  1981 => (x"3e",x"1c",x"00",x"00"),
  1982 => (x"00",x"00",x"41",x"63"),
  1983 => (x"63",x"41",x"00",x"00"),
  1984 => (x"00",x"00",x"1c",x"3e"),
  1985 => (x"1c",x"3e",x"2a",x"08"),
  1986 => (x"08",x"2a",x"3e",x"1c"),
  1987 => (x"3e",x"08",x"08",x"00"),
  1988 => (x"00",x"08",x"08",x"3e"),
  1989 => (x"e0",x"80",x"00",x"00"),
  1990 => (x"00",x"00",x"00",x"60"),
  1991 => (x"08",x"08",x"08",x"00"),
  1992 => (x"00",x"08",x"08",x"08"),
  1993 => (x"60",x"00",x"00",x"00"),
  1994 => (x"00",x"00",x"00",x"60"),
  1995 => (x"18",x"30",x"60",x"40"),
  1996 => (x"01",x"03",x"06",x"0c"),
  1997 => (x"59",x"7f",x"3e",x"00"),
  1998 => (x"00",x"3e",x"7f",x"4d"),
  1999 => (x"7f",x"06",x"04",x"00"),
  2000 => (x"00",x"00",x"00",x"7f"),
  2001 => (x"71",x"63",x"42",x"00"),
  2002 => (x"00",x"46",x"4f",x"59"),
  2003 => (x"49",x"63",x"22",x"00"),
  2004 => (x"00",x"36",x"7f",x"49"),
  2005 => (x"13",x"16",x"1c",x"18"),
  2006 => (x"00",x"10",x"7f",x"7f"),
  2007 => (x"45",x"67",x"27",x"00"),
  2008 => (x"00",x"39",x"7d",x"45"),
  2009 => (x"4b",x"7e",x"3c",x"00"),
  2010 => (x"00",x"30",x"79",x"49"),
  2011 => (x"71",x"01",x"01",x"00"),
  2012 => (x"00",x"07",x"0f",x"79"),
  2013 => (x"49",x"7f",x"36",x"00"),
  2014 => (x"00",x"36",x"7f",x"49"),
  2015 => (x"49",x"4f",x"06",x"00"),
  2016 => (x"00",x"1e",x"3f",x"69"),
  2017 => (x"66",x"00",x"00",x"00"),
  2018 => (x"00",x"00",x"00",x"66"),
  2019 => (x"e6",x"80",x"00",x"00"),
  2020 => (x"00",x"00",x"00",x"66"),
  2021 => (x"14",x"08",x"08",x"00"),
  2022 => (x"00",x"22",x"22",x"14"),
  2023 => (x"14",x"14",x"14",x"00"),
  2024 => (x"00",x"14",x"14",x"14"),
  2025 => (x"14",x"22",x"22",x"00"),
  2026 => (x"00",x"08",x"08",x"14"),
  2027 => (x"51",x"03",x"02",x"00"),
  2028 => (x"00",x"06",x"0f",x"59"),
  2029 => (x"5d",x"41",x"7f",x"3e"),
  2030 => (x"00",x"1e",x"1f",x"55"),
  2031 => (x"09",x"7f",x"7e",x"00"),
  2032 => (x"00",x"7e",x"7f",x"09"),
  2033 => (x"49",x"7f",x"7f",x"00"),
  2034 => (x"00",x"36",x"7f",x"49"),
  2035 => (x"63",x"3e",x"1c",x"00"),
  2036 => (x"00",x"41",x"41",x"41"),
  2037 => (x"41",x"7f",x"7f",x"00"),
  2038 => (x"00",x"1c",x"3e",x"63"),
  2039 => (x"49",x"7f",x"7f",x"00"),
  2040 => (x"00",x"41",x"41",x"49"),
  2041 => (x"09",x"7f",x"7f",x"00"),
  2042 => (x"00",x"01",x"01",x"09"),
  2043 => (x"41",x"7f",x"3e",x"00"),
  2044 => (x"00",x"7a",x"7b",x"49"),
  2045 => (x"08",x"7f",x"7f",x"00"),
  2046 => (x"00",x"7f",x"7f",x"08"),
  2047 => (x"7f",x"41",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

