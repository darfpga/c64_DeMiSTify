
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"00",x"41",x"7f"),
     1 => (x"40",x"60",x"20",x"00"),
     2 => (x"00",x"3f",x"7f",x"40"),
     3 => (x"1c",x"08",x"7f",x"7f"),
     4 => (x"00",x"41",x"63",x"36"),
     5 => (x"40",x"7f",x"7f",x"00"),
     6 => (x"00",x"40",x"40",x"40"),
     7 => (x"0c",x"06",x"7f",x"7f"),
     8 => (x"00",x"7f",x"7f",x"06"),
     9 => (x"0c",x"06",x"7f",x"7f"),
    10 => (x"00",x"7f",x"7f",x"18"),
    11 => (x"41",x"7f",x"3e",x"00"),
    12 => (x"00",x"3e",x"7f",x"41"),
    13 => (x"09",x"7f",x"7f",x"00"),
    14 => (x"00",x"06",x"0f",x"09"),
    15 => (x"61",x"41",x"7f",x"3e"),
    16 => (x"00",x"40",x"7e",x"7f"),
    17 => (x"09",x"7f",x"7f",x"00"),
    18 => (x"00",x"66",x"7f",x"19"),
    19 => (x"4d",x"6f",x"26",x"00"),
    20 => (x"00",x"32",x"7b",x"59"),
    21 => (x"7f",x"01",x"01",x"00"),
    22 => (x"00",x"01",x"01",x"7f"),
    23 => (x"40",x"7f",x"3f",x"00"),
    24 => (x"00",x"3f",x"7f",x"40"),
    25 => (x"70",x"3f",x"0f",x"00"),
    26 => (x"00",x"0f",x"3f",x"70"),
    27 => (x"18",x"30",x"7f",x"7f"),
    28 => (x"00",x"7f",x"7f",x"30"),
    29 => (x"1c",x"36",x"63",x"41"),
    30 => (x"41",x"63",x"36",x"1c"),
    31 => (x"7c",x"06",x"03",x"01"),
    32 => (x"01",x"03",x"06",x"7c"),
    33 => (x"4d",x"59",x"71",x"61"),
    34 => (x"00",x"41",x"43",x"47"),
    35 => (x"7f",x"7f",x"00",x"00"),
    36 => (x"00",x"00",x"41",x"41"),
    37 => (x"0c",x"06",x"03",x"01"),
    38 => (x"40",x"60",x"30",x"18"),
    39 => (x"41",x"41",x"00",x"00"),
    40 => (x"00",x"00",x"7f",x"7f"),
    41 => (x"03",x"06",x"0c",x"08"),
    42 => (x"00",x"08",x"0c",x"06"),
    43 => (x"80",x"80",x"80",x"80"),
    44 => (x"00",x"80",x"80",x"80"),
    45 => (x"03",x"00",x"00",x"00"),
    46 => (x"00",x"00",x"04",x"07"),
    47 => (x"54",x"74",x"20",x"00"),
    48 => (x"00",x"78",x"7c",x"54"),
    49 => (x"44",x"7f",x"7f",x"00"),
    50 => (x"00",x"38",x"7c",x"44"),
    51 => (x"44",x"7c",x"38",x"00"),
    52 => (x"00",x"00",x"44",x"44"),
    53 => (x"44",x"7c",x"38",x"00"),
    54 => (x"00",x"7f",x"7f",x"44"),
    55 => (x"54",x"7c",x"38",x"00"),
    56 => (x"00",x"18",x"5c",x"54"),
    57 => (x"7f",x"7e",x"04",x"00"),
    58 => (x"00",x"00",x"05",x"05"),
    59 => (x"a4",x"bc",x"18",x"00"),
    60 => (x"00",x"7c",x"fc",x"a4"),
    61 => (x"04",x"7f",x"7f",x"00"),
    62 => (x"00",x"78",x"7c",x"04"),
    63 => (x"3d",x"00",x"00",x"00"),
    64 => (x"00",x"00",x"40",x"7d"),
    65 => (x"80",x"80",x"80",x"00"),
    66 => (x"00",x"00",x"7d",x"fd"),
    67 => (x"10",x"7f",x"7f",x"00"),
    68 => (x"00",x"44",x"6c",x"38"),
    69 => (x"3f",x"00",x"00",x"00"),
    70 => (x"00",x"00",x"40",x"7f"),
    71 => (x"18",x"0c",x"7c",x"7c"),
    72 => (x"00",x"78",x"7c",x"0c"),
    73 => (x"04",x"7c",x"7c",x"00"),
    74 => (x"00",x"78",x"7c",x"04"),
    75 => (x"44",x"7c",x"38",x"00"),
    76 => (x"00",x"38",x"7c",x"44"),
    77 => (x"24",x"fc",x"fc",x"00"),
    78 => (x"00",x"18",x"3c",x"24"),
    79 => (x"24",x"3c",x"18",x"00"),
    80 => (x"00",x"fc",x"fc",x"24"),
    81 => (x"04",x"7c",x"7c",x"00"),
    82 => (x"00",x"08",x"0c",x"04"),
    83 => (x"54",x"5c",x"48",x"00"),
    84 => (x"00",x"20",x"74",x"54"),
    85 => (x"7f",x"3f",x"04",x"00"),
    86 => (x"00",x"00",x"44",x"44"),
    87 => (x"40",x"7c",x"3c",x"00"),
    88 => (x"00",x"7c",x"7c",x"40"),
    89 => (x"60",x"3c",x"1c",x"00"),
    90 => (x"00",x"1c",x"3c",x"60"),
    91 => (x"30",x"60",x"7c",x"3c"),
    92 => (x"00",x"3c",x"7c",x"60"),
    93 => (x"10",x"38",x"6c",x"44"),
    94 => (x"00",x"44",x"6c",x"38"),
    95 => (x"e0",x"bc",x"1c",x"00"),
    96 => (x"00",x"1c",x"3c",x"60"),
    97 => (x"74",x"64",x"44",x"00"),
    98 => (x"00",x"44",x"4c",x"5c"),
    99 => (x"3e",x"08",x"08",x"00"),
   100 => (x"00",x"41",x"41",x"77"),
   101 => (x"7f",x"00",x"00",x"00"),
   102 => (x"00",x"00",x"00",x"7f"),
   103 => (x"77",x"41",x"41",x"00"),
   104 => (x"00",x"08",x"08",x"3e"),
   105 => (x"03",x"01",x"01",x"02"),
   106 => (x"00",x"01",x"02",x"02"),
   107 => (x"7f",x"7f",x"7f",x"7f"),
   108 => (x"00",x"7f",x"7f",x"7f"),
   109 => (x"1c",x"1c",x"08",x"08"),
   110 => (x"7f",x"7f",x"3e",x"3e"),
   111 => (x"3e",x"3e",x"7f",x"7f"),
   112 => (x"08",x"08",x"1c",x"1c"),
   113 => (x"7c",x"18",x"10",x"00"),
   114 => (x"00",x"10",x"18",x"7c"),
   115 => (x"7c",x"30",x"10",x"00"),
   116 => (x"00",x"10",x"30",x"7c"),
   117 => (x"60",x"60",x"30",x"10"),
   118 => (x"00",x"06",x"1e",x"78"),
   119 => (x"18",x"3c",x"66",x"42"),
   120 => (x"00",x"42",x"66",x"3c"),
   121 => (x"c2",x"6a",x"38",x"78"),
   122 => (x"00",x"38",x"6c",x"c6"),
   123 => (x"60",x"00",x"00",x"60"),
   124 => (x"00",x"60",x"00",x"00"),
   125 => (x"5c",x"5b",x"5e",x"0e"),
   126 => (x"71",x"1e",x"0e",x"5d"),
   127 => (x"d9",x"f1",x"c2",x"4c"),
   128 => (x"4b",x"c0",x"4d",x"bf"),
   129 => (x"ab",x"74",x"1e",x"c0"),
   130 => (x"c4",x"87",x"c7",x"02"),
   131 => (x"78",x"c0",x"48",x"a6"),
   132 => (x"a6",x"c4",x"87",x"c5"),
   133 => (x"c4",x"78",x"c1",x"48"),
   134 => (x"49",x"73",x"1e",x"66"),
   135 => (x"c8",x"87",x"df",x"ee"),
   136 => (x"49",x"e0",x"c0",x"86"),
   137 => (x"c4",x"87",x"ef",x"ef"),
   138 => (x"49",x"6a",x"4a",x"a5"),
   139 => (x"f1",x"87",x"f0",x"f0"),
   140 => (x"85",x"cb",x"87",x"c6"),
   141 => (x"b7",x"c8",x"83",x"c1"),
   142 => (x"c7",x"ff",x"04",x"ab"),
   143 => (x"4d",x"26",x"26",x"87"),
   144 => (x"4b",x"26",x"4c",x"26"),
   145 => (x"71",x"1e",x"4f",x"26"),
   146 => (x"dd",x"f1",x"c2",x"4a"),
   147 => (x"dd",x"f1",x"c2",x"5a"),
   148 => (x"49",x"78",x"c7",x"48"),
   149 => (x"26",x"87",x"dd",x"fe"),
   150 => (x"1e",x"73",x"1e",x"4f"),
   151 => (x"b7",x"c0",x"4a",x"71"),
   152 => (x"87",x"d3",x"03",x"aa"),
   153 => (x"bf",x"f3",x"d6",x"c2"),
   154 => (x"c1",x"87",x"c4",x"05"),
   155 => (x"c0",x"87",x"c2",x"4b"),
   156 => (x"f7",x"d6",x"c2",x"4b"),
   157 => (x"c2",x"87",x"c4",x"5b"),
   158 => (x"c2",x"5a",x"f7",x"d6"),
   159 => (x"4a",x"bf",x"f3",x"d6"),
   160 => (x"c0",x"c1",x"9a",x"c1"),
   161 => (x"e8",x"ec",x"49",x"a2"),
   162 => (x"c2",x"48",x"fc",x"87"),
   163 => (x"78",x"bf",x"f3",x"d6"),
   164 => (x"1e",x"87",x"ef",x"fe"),
   165 => (x"66",x"c4",x"4a",x"71"),
   166 => (x"e6",x"49",x"72",x"1e"),
   167 => (x"26",x"26",x"87",x"e2"),
   168 => (x"d6",x"c2",x"1e",x"4f"),
   169 => (x"e3",x"49",x"bf",x"f3"),
   170 => (x"f1",x"c2",x"87",x"c4"),
   171 => (x"bf",x"e8",x"48",x"d1"),
   172 => (x"cd",x"f1",x"c2",x"78"),
   173 => (x"78",x"bf",x"ec",x"48"),
   174 => (x"bf",x"d1",x"f1",x"c2"),
   175 => (x"ff",x"c3",x"49",x"4a"),
   176 => (x"2a",x"b7",x"c8",x"99"),
   177 => (x"b0",x"71",x"48",x"72"),
   178 => (x"58",x"d9",x"f1",x"c2"),
   179 => (x"5e",x"0e",x"4f",x"26"),
   180 => (x"0e",x"5d",x"5c",x"5b"),
   181 => (x"c8",x"ff",x"4b",x"71"),
   182 => (x"cc",x"f1",x"c2",x"87"),
   183 => (x"73",x"50",x"c0",x"48"),
   184 => (x"87",x"ea",x"e2",x"49"),
   185 => (x"c2",x"4c",x"49",x"70"),
   186 => (x"49",x"ee",x"cb",x"9c"),
   187 => (x"70",x"87",x"cc",x"cb"),
   188 => (x"f1",x"c2",x"4d",x"49"),
   189 => (x"05",x"bf",x"97",x"cc"),
   190 => (x"d0",x"87",x"e2",x"c1"),
   191 => (x"f1",x"c2",x"49",x"66"),
   192 => (x"05",x"99",x"bf",x"d5"),
   193 => (x"66",x"d4",x"87",x"d6"),
   194 => (x"cd",x"f1",x"c2",x"49"),
   195 => (x"cb",x"05",x"99",x"bf"),
   196 => (x"e1",x"49",x"73",x"87"),
   197 => (x"98",x"70",x"87",x"f8"),
   198 => (x"87",x"c1",x"c1",x"02"),
   199 => (x"c0",x"fe",x"4c",x"c1"),
   200 => (x"ca",x"49",x"75",x"87"),
   201 => (x"98",x"70",x"87",x"e1"),
   202 => (x"c2",x"87",x"c6",x"02"),
   203 => (x"c1",x"48",x"cc",x"f1"),
   204 => (x"cc",x"f1",x"c2",x"50"),
   205 => (x"c0",x"05",x"bf",x"97"),
   206 => (x"f1",x"c2",x"87",x"e3"),
   207 => (x"d0",x"49",x"bf",x"d5"),
   208 => (x"ff",x"05",x"99",x"66"),
   209 => (x"f1",x"c2",x"87",x"d6"),
   210 => (x"d4",x"49",x"bf",x"cd"),
   211 => (x"ff",x"05",x"99",x"66"),
   212 => (x"49",x"73",x"87",x"ca"),
   213 => (x"70",x"87",x"f7",x"e0"),
   214 => (x"ff",x"fe",x"05",x"98"),
   215 => (x"fb",x"48",x"74",x"87"),
   216 => (x"5e",x"0e",x"87",x"dc"),
   217 => (x"0e",x"5d",x"5c",x"5b"),
   218 => (x"4d",x"c0",x"86",x"f4"),
   219 => (x"7e",x"bf",x"ec",x"4c"),
   220 => (x"c2",x"48",x"a6",x"c4"),
   221 => (x"78",x"bf",x"d9",x"f1"),
   222 => (x"1e",x"c0",x"1e",x"c1"),
   223 => (x"cd",x"fd",x"49",x"c7"),
   224 => (x"70",x"86",x"c8",x"87"),
   225 => (x"87",x"ce",x"02",x"98"),
   226 => (x"cc",x"fb",x"49",x"ff"),
   227 => (x"49",x"da",x"c1",x"87"),
   228 => (x"87",x"fa",x"df",x"ff"),
   229 => (x"f1",x"c2",x"4d",x"c1"),
   230 => (x"02",x"bf",x"97",x"cc"),
   231 => (x"c4",x"d0",x"87",x"c3"),
   232 => (x"d1",x"f1",x"c2",x"87"),
   233 => (x"d6",x"c2",x"4b",x"bf"),
   234 => (x"c0",x"05",x"bf",x"f3"),
   235 => (x"fd",x"c3",x"87",x"eb"),
   236 => (x"d9",x"df",x"ff",x"49"),
   237 => (x"49",x"fa",x"c3",x"87"),
   238 => (x"87",x"d2",x"df",x"ff"),
   239 => (x"ff",x"c3",x"49",x"73"),
   240 => (x"c0",x"1e",x"71",x"99"),
   241 => (x"87",x"cb",x"fb",x"49"),
   242 => (x"b7",x"c8",x"49",x"73"),
   243 => (x"c1",x"1e",x"71",x"29"),
   244 => (x"87",x"ff",x"fa",x"49"),
   245 => (x"c0",x"c6",x"86",x"c8"),
   246 => (x"d5",x"f1",x"c2",x"87"),
   247 => (x"02",x"9b",x"4b",x"bf"),
   248 => (x"d6",x"c2",x"87",x"dd"),
   249 => (x"c7",x"49",x"bf",x"ef"),
   250 => (x"98",x"70",x"87",x"dd"),
   251 => (x"c0",x"87",x"c4",x"05"),
   252 => (x"c2",x"87",x"d2",x"4b"),
   253 => (x"c2",x"c7",x"49",x"e0"),
   254 => (x"f3",x"d6",x"c2",x"87"),
   255 => (x"c2",x"87",x"c6",x"58"),
   256 => (x"c0",x"48",x"ef",x"d6"),
   257 => (x"c2",x"49",x"73",x"78"),
   258 => (x"87",x"ce",x"05",x"99"),
   259 => (x"ff",x"49",x"eb",x"c3"),
   260 => (x"70",x"87",x"fb",x"dd"),
   261 => (x"02",x"99",x"c2",x"49"),
   262 => (x"4c",x"fb",x"87",x"c2"),
   263 => (x"99",x"c1",x"49",x"73"),
   264 => (x"c3",x"87",x"ce",x"05"),
   265 => (x"dd",x"ff",x"49",x"f4"),
   266 => (x"49",x"70",x"87",x"e4"),
   267 => (x"c2",x"02",x"99",x"c2"),
   268 => (x"73",x"4c",x"fa",x"87"),
   269 => (x"05",x"99",x"c8",x"49"),
   270 => (x"f5",x"c3",x"87",x"ce"),
   271 => (x"cd",x"dd",x"ff",x"49"),
   272 => (x"c2",x"49",x"70",x"87"),
   273 => (x"87",x"d5",x"02",x"99"),
   274 => (x"bf",x"dd",x"f1",x"c2"),
   275 => (x"48",x"87",x"ca",x"02"),
   276 => (x"f1",x"c2",x"88",x"c1"),
   277 => (x"c2",x"c0",x"58",x"e1"),
   278 => (x"c1",x"4c",x"ff",x"87"),
   279 => (x"c4",x"49",x"73",x"4d"),
   280 => (x"87",x"ce",x"05",x"99"),
   281 => (x"ff",x"49",x"f2",x"c3"),
   282 => (x"70",x"87",x"e3",x"dc"),
   283 => (x"02",x"99",x"c2",x"49"),
   284 => (x"f1",x"c2",x"87",x"dc"),
   285 => (x"48",x"7e",x"bf",x"dd"),
   286 => (x"03",x"a8",x"b7",x"c7"),
   287 => (x"6e",x"87",x"cb",x"c0"),
   288 => (x"c2",x"80",x"c1",x"48"),
   289 => (x"c0",x"58",x"e1",x"f1"),
   290 => (x"4c",x"fe",x"87",x"c2"),
   291 => (x"fd",x"c3",x"4d",x"c1"),
   292 => (x"f9",x"db",x"ff",x"49"),
   293 => (x"c2",x"49",x"70",x"87"),
   294 => (x"87",x"d5",x"02",x"99"),
   295 => (x"bf",x"dd",x"f1",x"c2"),
   296 => (x"87",x"c9",x"c0",x"02"),
   297 => (x"48",x"dd",x"f1",x"c2"),
   298 => (x"c2",x"c0",x"78",x"c0"),
   299 => (x"c1",x"4c",x"fd",x"87"),
   300 => (x"49",x"fa",x"c3",x"4d"),
   301 => (x"87",x"d6",x"db",x"ff"),
   302 => (x"99",x"c2",x"49",x"70"),
   303 => (x"87",x"d9",x"c0",x"02"),
   304 => (x"bf",x"dd",x"f1",x"c2"),
   305 => (x"a8",x"b7",x"c7",x"48"),
   306 => (x"87",x"c9",x"c0",x"03"),
   307 => (x"48",x"dd",x"f1",x"c2"),
   308 => (x"c2",x"c0",x"78",x"c7"),
   309 => (x"c1",x"4c",x"fc",x"87"),
   310 => (x"ac",x"b7",x"c0",x"4d"),
   311 => (x"87",x"d1",x"c0",x"03"),
   312 => (x"c1",x"4a",x"66",x"c4"),
   313 => (x"02",x"6a",x"82",x"d8"),
   314 => (x"6a",x"87",x"c6",x"c0"),
   315 => (x"73",x"49",x"74",x"4b"),
   316 => (x"c3",x"1e",x"c0",x"0f"),
   317 => (x"da",x"c1",x"1e",x"f0"),
   318 => (x"87",x"d2",x"f7",x"49"),
   319 => (x"98",x"70",x"86",x"c8"),
   320 => (x"87",x"e2",x"c0",x"02"),
   321 => (x"c2",x"48",x"a6",x"c8"),
   322 => (x"78",x"bf",x"dd",x"f1"),
   323 => (x"cb",x"49",x"66",x"c8"),
   324 => (x"48",x"66",x"c4",x"91"),
   325 => (x"7e",x"70",x"80",x"71"),
   326 => (x"c0",x"02",x"bf",x"6e"),
   327 => (x"bf",x"6e",x"87",x"c8"),
   328 => (x"49",x"66",x"c8",x"4b"),
   329 => (x"9d",x"75",x"0f",x"73"),
   330 => (x"87",x"c8",x"c0",x"02"),
   331 => (x"bf",x"dd",x"f1",x"c2"),
   332 => (x"87",x"c0",x"f3",x"49"),
   333 => (x"bf",x"f7",x"d6",x"c2"),
   334 => (x"87",x"dd",x"c0",x"02"),
   335 => (x"87",x"c7",x"c2",x"49"),
   336 => (x"c0",x"02",x"98",x"70"),
   337 => (x"f1",x"c2",x"87",x"d3"),
   338 => (x"f2",x"49",x"bf",x"dd"),
   339 => (x"49",x"c0",x"87",x"e6"),
   340 => (x"c2",x"87",x"c6",x"f4"),
   341 => (x"c0",x"48",x"f7",x"d6"),
   342 => (x"f3",x"8e",x"f4",x"78"),
   343 => (x"5e",x"0e",x"87",x"e0"),
   344 => (x"0e",x"5d",x"5c",x"5b"),
   345 => (x"c2",x"4c",x"71",x"1e"),
   346 => (x"49",x"bf",x"d9",x"f1"),
   347 => (x"4d",x"a1",x"cd",x"c1"),
   348 => (x"69",x"81",x"d1",x"c1"),
   349 => (x"02",x"9c",x"74",x"7e"),
   350 => (x"a5",x"c4",x"87",x"cf"),
   351 => (x"c2",x"7b",x"74",x"4b"),
   352 => (x"49",x"bf",x"d9",x"f1"),
   353 => (x"6e",x"87",x"ff",x"f2"),
   354 => (x"05",x"9c",x"74",x"7b"),
   355 => (x"4b",x"c0",x"87",x"c4"),
   356 => (x"4b",x"c1",x"87",x"c2"),
   357 => (x"c0",x"f3",x"49",x"73"),
   358 => (x"02",x"66",x"d4",x"87"),
   359 => (x"da",x"49",x"87",x"c7"),
   360 => (x"c2",x"4a",x"70",x"87"),
   361 => (x"c2",x"4a",x"c0",x"87"),
   362 => (x"26",x"5a",x"fb",x"d6"),
   363 => (x"00",x"87",x"cf",x"f2"),
   364 => (x"00",x"00",x"00",x"00"),
   365 => (x"00",x"00",x"00",x"00"),
   366 => (x"1e",x"00",x"00",x"00"),
   367 => (x"c8",x"ff",x"4a",x"71"),
   368 => (x"a1",x"72",x"49",x"bf"),
   369 => (x"1e",x"4f",x"26",x"48"),
   370 => (x"89",x"bf",x"c8",x"ff"),
   371 => (x"c0",x"c0",x"c0",x"fe"),
   372 => (x"01",x"a9",x"c0",x"c0"),
   373 => (x"4a",x"c0",x"87",x"c4"),
   374 => (x"4a",x"c1",x"87",x"c2"),
   375 => (x"4f",x"26",x"48",x"72"),
   376 => (x"5c",x"5b",x"5e",x"0e"),
   377 => (x"4b",x"71",x"0e",x"5d"),
   378 => (x"d0",x"4c",x"d4",x"ff"),
   379 => (x"78",x"c0",x"48",x"66"),
   380 => (x"d8",x"ff",x"49",x"d6"),
   381 => (x"ff",x"c3",x"87",x"d0"),
   382 => (x"c3",x"49",x"6c",x"7c"),
   383 => (x"4d",x"71",x"99",x"ff"),
   384 => (x"99",x"f0",x"c3",x"49"),
   385 => (x"05",x"a9",x"e0",x"c1"),
   386 => (x"ff",x"c3",x"87",x"cb"),
   387 => (x"c3",x"48",x"6c",x"7c"),
   388 => (x"08",x"66",x"d0",x"98"),
   389 => (x"7c",x"ff",x"c3",x"78"),
   390 => (x"c8",x"49",x"4a",x"6c"),
   391 => (x"7c",x"ff",x"c3",x"31"),
   392 => (x"b2",x"71",x"4a",x"6c"),
   393 => (x"31",x"c8",x"49",x"72"),
   394 => (x"6c",x"7c",x"ff",x"c3"),
   395 => (x"72",x"b2",x"71",x"4a"),
   396 => (x"c3",x"31",x"c8",x"49"),
   397 => (x"4a",x"6c",x"7c",x"ff"),
   398 => (x"d0",x"ff",x"b2",x"71"),
   399 => (x"78",x"e0",x"c0",x"48"),
   400 => (x"c2",x"02",x"9b",x"73"),
   401 => (x"75",x"7b",x"72",x"87"),
   402 => (x"26",x"4d",x"26",x"48"),
   403 => (x"26",x"4b",x"26",x"4c"),
   404 => (x"4f",x"26",x"1e",x"4f"),
   405 => (x"5c",x"5b",x"5e",x"0e"),
   406 => (x"76",x"86",x"f8",x"0e"),
   407 => (x"49",x"a6",x"c8",x"1e"),
   408 => (x"c4",x"87",x"fd",x"fd"),
   409 => (x"6e",x"4b",x"70",x"86"),
   410 => (x"03",x"a8",x"c2",x"48"),
   411 => (x"73",x"87",x"f0",x"c2"),
   412 => (x"9a",x"f0",x"c3",x"4a"),
   413 => (x"02",x"aa",x"d0",x"c1"),
   414 => (x"e0",x"c1",x"87",x"c7"),
   415 => (x"de",x"c2",x"05",x"aa"),
   416 => (x"c8",x"49",x"73",x"87"),
   417 => (x"87",x"c3",x"02",x"99"),
   418 => (x"73",x"87",x"c6",x"ff"),
   419 => (x"c2",x"9c",x"c3",x"4c"),
   420 => (x"c2",x"c1",x"05",x"ac"),
   421 => (x"49",x"66",x"c4",x"87"),
   422 => (x"1e",x"71",x"31",x"c9"),
   423 => (x"d4",x"4a",x"66",x"c4"),
   424 => (x"e1",x"f1",x"c2",x"92"),
   425 => (x"fe",x"81",x"72",x"49"),
   426 => (x"d8",x"87",x"e7",x"cc"),
   427 => (x"d5",x"d5",x"ff",x"49"),
   428 => (x"1e",x"c0",x"c8",x"87"),
   429 => (x"49",x"fa",x"df",x"c2"),
   430 => (x"87",x"e3",x"e8",x"fd"),
   431 => (x"c0",x"48",x"d0",x"ff"),
   432 => (x"df",x"c2",x"78",x"e0"),
   433 => (x"66",x"cc",x"1e",x"fa"),
   434 => (x"c2",x"92",x"d4",x"4a"),
   435 => (x"72",x"49",x"e1",x"f1"),
   436 => (x"ee",x"ca",x"fe",x"81"),
   437 => (x"c1",x"86",x"cc",x"87"),
   438 => (x"c2",x"c1",x"05",x"ac"),
   439 => (x"49",x"66",x"c4",x"87"),
   440 => (x"1e",x"71",x"31",x"c9"),
   441 => (x"d4",x"4a",x"66",x"c4"),
   442 => (x"e1",x"f1",x"c2",x"92"),
   443 => (x"fe",x"81",x"72",x"49"),
   444 => (x"c2",x"87",x"df",x"cb"),
   445 => (x"c8",x"1e",x"fa",x"df"),
   446 => (x"92",x"d4",x"4a",x"66"),
   447 => (x"49",x"e1",x"f1",x"c2"),
   448 => (x"c8",x"fe",x"81",x"72"),
   449 => (x"49",x"d7",x"87",x"ee"),
   450 => (x"87",x"fa",x"d3",x"ff"),
   451 => (x"c2",x"1e",x"c0",x"c8"),
   452 => (x"fd",x"49",x"fa",x"df"),
   453 => (x"cc",x"87",x"e1",x"e6"),
   454 => (x"48",x"d0",x"ff",x"86"),
   455 => (x"f8",x"78",x"e0",x"c0"),
   456 => (x"87",x"e7",x"fc",x"8e"),
   457 => (x"5c",x"5b",x"5e",x"0e"),
   458 => (x"71",x"1e",x"0e",x"5d"),
   459 => (x"4c",x"d4",x"ff",x"4d"),
   460 => (x"48",x"7e",x"66",x"d4"),
   461 => (x"06",x"a8",x"b7",x"c3"),
   462 => (x"48",x"c0",x"87",x"c5"),
   463 => (x"75",x"87",x"e2",x"c1"),
   464 => (x"f2",x"d9",x"fe",x"49"),
   465 => (x"c4",x"1e",x"75",x"87"),
   466 => (x"93",x"d4",x"4b",x"66"),
   467 => (x"83",x"e1",x"f1",x"c2"),
   468 => (x"c2",x"fe",x"49",x"73"),
   469 => (x"83",x"c8",x"87",x"eb"),
   470 => (x"d0",x"ff",x"4b",x"6b"),
   471 => (x"78",x"e1",x"c8",x"48"),
   472 => (x"49",x"73",x"7c",x"dd"),
   473 => (x"71",x"99",x"ff",x"c3"),
   474 => (x"c8",x"49",x"73",x"7c"),
   475 => (x"ff",x"c3",x"29",x"b7"),
   476 => (x"73",x"7c",x"71",x"99"),
   477 => (x"29",x"b7",x"d0",x"49"),
   478 => (x"71",x"99",x"ff",x"c3"),
   479 => (x"d8",x"49",x"73",x"7c"),
   480 => (x"7c",x"71",x"29",x"b7"),
   481 => (x"7c",x"7c",x"7c",x"c0"),
   482 => (x"7c",x"7c",x"7c",x"7c"),
   483 => (x"7c",x"7c",x"7c",x"7c"),
   484 => (x"78",x"e0",x"c0",x"7c"),
   485 => (x"dc",x"1e",x"66",x"c4"),
   486 => (x"ce",x"d2",x"ff",x"49"),
   487 => (x"73",x"86",x"c8",x"87"),
   488 => (x"e4",x"fa",x"26",x"48"),
   489 => (x"df",x"c2",x"1e",x"87"),
   490 => (x"c1",x"49",x"bf",x"ce"),
   491 => (x"d2",x"df",x"c2",x"b9"),
   492 => (x"48",x"d4",x"ff",x"59"),
   493 => (x"ff",x"78",x"ff",x"c3"),
   494 => (x"e1",x"c0",x"48",x"d0"),
   495 => (x"48",x"d4",x"ff",x"78"),
   496 => (x"31",x"c4",x"78",x"c1"),
   497 => (x"d0",x"ff",x"78",x"71"),
   498 => (x"78",x"e0",x"c0",x"48"),
   499 => (x"00",x"00",x"4f",x"26"),
   500 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

